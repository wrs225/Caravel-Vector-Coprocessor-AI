magic
tech sky130A
magscale 1 2
timestamp 1692295508
<< obsli1 >>
rect 1104 2159 243156 183345
<< obsm1 >>
rect 14 892 243418 185088
<< metal2 >>
rect 5814 185138 5870 185938
rect 12898 185138 12954 185938
rect 19338 185138 19394 185938
rect 25778 185138 25834 185938
rect 32218 185138 32274 185938
rect 38658 185138 38714 185938
rect 45098 185138 45154 185938
rect 51538 185138 51594 185938
rect 58622 185138 58678 185938
rect 65062 185138 65118 185938
rect 71502 185138 71558 185938
rect 77942 185138 77998 185938
rect 84382 185138 84438 185938
rect 90822 185138 90878 185938
rect 97262 185138 97318 185938
rect 103702 185138 103758 185938
rect 110786 185138 110842 185938
rect 117226 185138 117282 185938
rect 123666 185138 123722 185938
rect 130106 185138 130162 185938
rect 136546 185138 136602 185938
rect 142986 185138 143042 185938
rect 149426 185138 149482 185938
rect 156510 185138 156566 185938
rect 162950 185138 163006 185938
rect 169390 185138 169446 185938
rect 175830 185138 175886 185938
rect 182270 185138 182326 185938
rect 188710 185138 188766 185938
rect 195150 185138 195206 185938
rect 202234 185138 202290 185938
rect 208674 185138 208730 185938
rect 215114 185138 215170 185938
rect 221554 185138 221610 185938
rect 227994 185138 228050 185938
rect 234434 185138 234490 185938
rect 240874 185138 240930 185938
rect 18 0 74 800
rect 6458 0 6514 800
rect 12898 0 12954 800
rect 19338 0 19394 800
rect 25778 0 25834 800
rect 32218 0 32274 800
rect 38658 0 38714 800
rect 45098 0 45154 800
rect 52182 0 52238 800
rect 58622 0 58678 800
rect 65062 0 65118 800
rect 71502 0 71558 800
rect 77942 0 77998 800
rect 84382 0 84438 800
rect 90822 0 90878 800
rect 97906 0 97962 800
rect 104346 0 104402 800
rect 110786 0 110842 800
rect 117226 0 117282 800
rect 123666 0 123722 800
rect 130106 0 130162 800
rect 136546 0 136602 800
rect 143630 0 143686 800
rect 150070 0 150126 800
rect 156510 0 156566 800
rect 162950 0 163006 800
rect 169390 0 169446 800
rect 175830 0 175886 800
rect 182270 0 182326 800
rect 189354 0 189410 800
rect 195794 0 195850 800
rect 202234 0 202290 800
rect 208674 0 208730 800
rect 215114 0 215170 800
rect 221554 0 221610 800
rect 227994 0 228050 800
rect 235078 0 235134 800
rect 241518 0 241574 800
<< obsm2 >>
rect 20 185082 5758 185745
rect 5926 185082 12842 185745
rect 13010 185082 19282 185745
rect 19450 185082 25722 185745
rect 25890 185082 32162 185745
rect 32330 185082 38602 185745
rect 38770 185082 45042 185745
rect 45210 185082 51482 185745
rect 51650 185082 58566 185745
rect 58734 185082 65006 185745
rect 65174 185082 71446 185745
rect 71614 185082 77886 185745
rect 78054 185082 84326 185745
rect 84494 185082 90766 185745
rect 90934 185082 97206 185745
rect 97374 185082 103646 185745
rect 103814 185082 110730 185745
rect 110898 185082 117170 185745
rect 117338 185082 123610 185745
rect 123778 185082 130050 185745
rect 130218 185082 136490 185745
rect 136658 185082 142930 185745
rect 143098 185082 149370 185745
rect 149538 185082 156454 185745
rect 156622 185082 162894 185745
rect 163062 185082 169334 185745
rect 169502 185082 175774 185745
rect 175942 185082 182214 185745
rect 182382 185082 188654 185745
rect 188822 185082 195094 185745
rect 195262 185082 202178 185745
rect 202346 185082 208618 185745
rect 208786 185082 215058 185745
rect 215226 185082 221498 185745
rect 221666 185082 227938 185745
rect 228106 185082 234378 185745
rect 234546 185082 240818 185745
rect 240986 185082 243414 185745
rect 20 856 243414 185082
rect 130 734 6402 856
rect 6570 734 12842 856
rect 13010 734 19282 856
rect 19450 734 25722 856
rect 25890 734 32162 856
rect 32330 734 38602 856
rect 38770 734 45042 856
rect 45210 734 52126 856
rect 52294 734 58566 856
rect 58734 734 65006 856
rect 65174 734 71446 856
rect 71614 734 77886 856
rect 78054 734 84326 856
rect 84494 734 90766 856
rect 90934 734 97850 856
rect 98018 734 104290 856
rect 104458 734 110730 856
rect 110898 734 117170 856
rect 117338 734 123610 856
rect 123778 734 130050 856
rect 130218 734 136490 856
rect 136658 734 143574 856
rect 143742 734 150014 856
rect 150182 734 156454 856
rect 156622 734 162894 856
rect 163062 734 169334 856
rect 169502 734 175774 856
rect 175942 734 182214 856
rect 182382 734 189298 856
rect 189466 734 195738 856
rect 195906 734 202178 856
rect 202346 734 208618 856
rect 208786 734 215058 856
rect 215226 734 221498 856
rect 221666 734 227938 856
rect 228106 734 235022 856
rect 235190 734 241462 856
rect 241630 734 243414 856
<< metal3 >>
rect 0 185648 800 185768
rect 243523 182248 244323 182368
rect 0 178848 800 178968
rect 243523 175448 244323 175568
rect 0 172048 800 172168
rect 243523 168648 244323 168768
rect 0 165248 800 165368
rect 243523 161848 244323 161968
rect 0 158448 800 158568
rect 243523 155048 244323 155168
rect 0 151648 800 151768
rect 243523 148248 244323 148368
rect 0 144168 800 144288
rect 243523 141448 244323 141568
rect 0 137368 800 137488
rect 243523 133968 244323 134088
rect 0 130568 800 130688
rect 243523 127168 244323 127288
rect 0 123768 800 123888
rect 243523 120368 244323 120488
rect 0 116968 800 117088
rect 243523 113568 244323 113688
rect 0 110168 800 110288
rect 243523 106768 244323 106888
rect 0 103368 800 103488
rect 243523 99968 244323 100088
rect 0 95888 800 96008
rect 243523 93168 244323 93288
rect 0 89088 800 89208
rect 243523 85688 244323 85808
rect 0 82288 800 82408
rect 243523 78888 244323 79008
rect 0 75488 800 75608
rect 243523 72088 244323 72208
rect 0 68688 800 68808
rect 243523 65288 244323 65408
rect 0 61888 800 62008
rect 243523 58488 244323 58608
rect 0 55088 800 55208
rect 243523 51688 244323 51808
rect 0 47608 800 47728
rect 243523 44888 244323 45008
rect 0 40808 800 40928
rect 243523 38088 244323 38208
rect 0 34008 800 34128
rect 243523 30608 244323 30728
rect 0 27208 800 27328
rect 243523 23808 244323 23928
rect 0 20408 800 20528
rect 243523 17008 244323 17128
rect 0 13608 800 13728
rect 243523 10208 244323 10328
rect 0 6808 800 6928
rect 243523 3408 244323 3528
<< obsm3 >>
rect 880 185568 243523 185741
rect 800 182448 243523 185568
rect 800 182168 243443 182448
rect 800 179048 243523 182168
rect 880 178768 243523 179048
rect 800 175648 243523 178768
rect 800 175368 243443 175648
rect 800 172248 243523 175368
rect 880 171968 243523 172248
rect 800 168848 243523 171968
rect 800 168568 243443 168848
rect 800 165448 243523 168568
rect 880 165168 243523 165448
rect 800 162048 243523 165168
rect 800 161768 243443 162048
rect 800 158648 243523 161768
rect 880 158368 243523 158648
rect 800 155248 243523 158368
rect 800 154968 243443 155248
rect 800 151848 243523 154968
rect 880 151568 243523 151848
rect 800 148448 243523 151568
rect 800 148168 243443 148448
rect 800 144368 243523 148168
rect 880 144088 243523 144368
rect 800 141648 243523 144088
rect 800 141368 243443 141648
rect 800 137568 243523 141368
rect 880 137288 243523 137568
rect 800 134168 243523 137288
rect 800 133888 243443 134168
rect 800 130768 243523 133888
rect 880 130488 243523 130768
rect 800 127368 243523 130488
rect 800 127088 243443 127368
rect 800 123968 243523 127088
rect 880 123688 243523 123968
rect 800 120568 243523 123688
rect 800 120288 243443 120568
rect 800 117168 243523 120288
rect 880 116888 243523 117168
rect 800 113768 243523 116888
rect 800 113488 243443 113768
rect 800 110368 243523 113488
rect 880 110088 243523 110368
rect 800 106968 243523 110088
rect 800 106688 243443 106968
rect 800 103568 243523 106688
rect 880 103288 243523 103568
rect 800 100168 243523 103288
rect 800 99888 243443 100168
rect 800 96088 243523 99888
rect 880 95808 243523 96088
rect 800 93368 243523 95808
rect 800 93088 243443 93368
rect 800 89288 243523 93088
rect 880 89008 243523 89288
rect 800 85888 243523 89008
rect 800 85608 243443 85888
rect 800 82488 243523 85608
rect 880 82208 243523 82488
rect 800 79088 243523 82208
rect 800 78808 243443 79088
rect 800 75688 243523 78808
rect 880 75408 243523 75688
rect 800 72288 243523 75408
rect 800 72008 243443 72288
rect 800 68888 243523 72008
rect 880 68608 243523 68888
rect 800 65488 243523 68608
rect 800 65208 243443 65488
rect 800 62088 243523 65208
rect 880 61808 243523 62088
rect 800 58688 243523 61808
rect 800 58408 243443 58688
rect 800 55288 243523 58408
rect 880 55008 243523 55288
rect 800 51888 243523 55008
rect 800 51608 243443 51888
rect 800 47808 243523 51608
rect 880 47528 243523 47808
rect 800 45088 243523 47528
rect 800 44808 243443 45088
rect 800 41008 243523 44808
rect 880 40728 243523 41008
rect 800 38288 243523 40728
rect 800 38008 243443 38288
rect 800 34208 243523 38008
rect 880 33928 243523 34208
rect 800 30808 243523 33928
rect 800 30528 243443 30808
rect 800 27408 243523 30528
rect 880 27128 243523 27408
rect 800 24008 243523 27128
rect 800 23728 243443 24008
rect 800 20608 243523 23728
rect 880 20328 243523 20608
rect 800 17208 243523 20328
rect 800 16928 243443 17208
rect 800 13808 243523 16928
rect 880 13528 243523 13808
rect 800 10408 243523 13528
rect 800 10128 243443 10408
rect 800 7008 243523 10128
rect 880 6728 243523 7008
rect 800 3608 243523 6728
rect 800 3328 243443 3608
rect 800 1531 243523 3328
<< metal4 >>
rect 4208 2128 4528 183376
rect 19568 2128 19888 183376
rect 34928 2128 35248 183376
rect 50288 2128 50608 183376
rect 65648 2128 65968 183376
rect 81008 2128 81328 183376
rect 96368 2128 96688 183376
rect 111728 2128 112048 183376
rect 127088 2128 127408 183376
rect 142448 2128 142768 183376
rect 157808 2128 158128 183376
rect 173168 2128 173488 183376
rect 188528 2128 188848 183376
rect 203888 2128 204208 183376
rect 219248 2128 219568 183376
rect 234608 2128 234928 183376
<< obsm4 >>
rect 4843 2048 19488 183157
rect 19968 2048 34848 183157
rect 35328 2048 50208 183157
rect 50688 2048 65568 183157
rect 66048 2048 80928 183157
rect 81408 2048 96288 183157
rect 96768 2048 111648 183157
rect 112128 2048 127008 183157
rect 127488 2048 142368 183157
rect 142848 2048 157728 183157
rect 158208 2048 173088 183157
rect 173568 2048 188448 183157
rect 188928 2048 203808 183157
rect 204288 2048 219168 183157
rect 219648 2048 234528 183157
rect 235008 2048 239509 183157
rect 4843 1531 239509 2048
<< labels >>
rlabel metal3 s 0 185648 800 185768 6 clk
port 1 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 rAddr1_1[0]
port 2 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 rAddr1_1[1]
port 3 nsew signal input
rlabel metal2 s 123666 185138 123722 185938 6 rAddr1_1[2]
port 4 nsew signal input
rlabel metal3 s 243523 182248 244323 182368 6 rAddr1_1[3]
port 5 nsew signal input
rlabel metal3 s 0 172048 800 172168 6 rAddr1_1[4]
port 6 nsew signal input
rlabel metal2 s 221554 185138 221610 185938 6 rAddr1_2[0]
port 7 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 rAddr1_2[1]
port 8 nsew signal input
rlabel metal2 s 65062 185138 65118 185938 6 rAddr1_2[2]
port 9 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 rAddr1_2[3]
port 10 nsew signal input
rlabel metal2 s 208674 185138 208730 185938 6 rAddr1_2[4]
port 11 nsew signal input
rlabel metal3 s 243523 51688 244323 51808 6 rAddr2_1[0]
port 12 nsew signal input
rlabel metal2 s 215114 185138 215170 185938 6 rAddr2_1[1]
port 13 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 rAddr2_1[2]
port 14 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 rAddr2_1[3]
port 15 nsew signal input
rlabel metal2 s 117226 185138 117282 185938 6 rAddr2_1[4]
port 16 nsew signal input
rlabel metal3 s 243523 44888 244323 45008 6 rAddr2_2[0]
port 17 nsew signal input
rlabel metal2 s 130106 185138 130162 185938 6 rAddr2_2[1]
port 18 nsew signal input
rlabel metal3 s 243523 127168 244323 127288 6 rAddr2_2[2]
port 19 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 rAddr2_2[3]
port 20 nsew signal input
rlabel metal3 s 243523 93168 244323 93288 6 rAddr2_2[4]
port 21 nsew signal input
rlabel metal3 s 243523 85688 244323 85808 6 rData1[0]
port 22 nsew signal output
rlabel metal2 s 77942 185138 77998 185938 6 rData1[10]
port 23 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 rData1[11]
port 24 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 rData1[12]
port 25 nsew signal output
rlabel metal3 s 243523 99968 244323 100088 6 rData1[13]
port 26 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 rData1[14]
port 27 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 rData1[15]
port 28 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 rData1[16]
port 29 nsew signal output
rlabel metal3 s 243523 120368 244323 120488 6 rData1[17]
port 30 nsew signal output
rlabel metal2 s 162950 185138 163006 185938 6 rData1[18]
port 31 nsew signal output
rlabel metal2 s 208674 0 208730 800 6 rData1[19]
port 32 nsew signal output
rlabel metal2 s 51538 185138 51594 185938 6 rData1[1]
port 33 nsew signal output
rlabel metal3 s 243523 30608 244323 30728 6 rData1[20]
port 34 nsew signal output
rlabel metal2 s 25778 185138 25834 185938 6 rData1[21]
port 35 nsew signal output
rlabel metal3 s 0 165248 800 165368 6 rData1[22]
port 36 nsew signal output
rlabel metal2 s 234434 185138 234490 185938 6 rData1[23]
port 37 nsew signal output
rlabel metal2 s 182270 0 182326 800 6 rData1[24]
port 38 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 rData1[25]
port 39 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 rData1[26]
port 40 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 rData1[27]
port 41 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 rData1[28]
port 42 nsew signal output
rlabel metal3 s 243523 10208 244323 10328 6 rData1[29]
port 43 nsew signal output
rlabel metal2 s 149426 185138 149482 185938 6 rData1[2]
port 44 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 rData1[30]
port 45 nsew signal output
rlabel metal2 s 182270 185138 182326 185938 6 rData1[31]
port 46 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 rData1[3]
port 47 nsew signal output
rlabel metal2 s 240874 185138 240930 185938 6 rData1[4]
port 48 nsew signal output
rlabel metal2 s 90822 185138 90878 185938 6 rData1[5]
port 49 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 rData1[6]
port 50 nsew signal output
rlabel metal3 s 243523 133968 244323 134088 6 rData1[7]
port 51 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 rData1[8]
port 52 nsew signal output
rlabel metal2 s 142986 185138 143042 185938 6 rData1[9]
port 53 nsew signal output
rlabel metal2 s 103702 185138 103758 185938 6 rData2[0]
port 54 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 rData2[10]
port 55 nsew signal output
rlabel metal3 s 243523 175448 244323 175568 6 rData2[11]
port 56 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 rData2[12]
port 57 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 rData2[13]
port 58 nsew signal output
rlabel metal2 s 84382 185138 84438 185938 6 rData2[14]
port 59 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 rData2[15]
port 60 nsew signal output
rlabel metal3 s 243523 161848 244323 161968 6 rData2[16]
port 61 nsew signal output
rlabel metal2 s 45098 185138 45154 185938 6 rData2[17]
port 62 nsew signal output
rlabel metal3 s 243523 148248 244323 148368 6 rData2[18]
port 63 nsew signal output
rlabel metal2 s 58622 185138 58678 185938 6 rData2[19]
port 64 nsew signal output
rlabel metal2 s 110786 185138 110842 185938 6 rData2[1]
port 65 nsew signal output
rlabel metal2 s 175830 185138 175886 185938 6 rData2[20]
port 66 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 rData2[21]
port 67 nsew signal output
rlabel metal3 s 243523 58488 244323 58608 6 rData2[22]
port 68 nsew signal output
rlabel metal3 s 243523 23808 244323 23928 6 rData2[23]
port 69 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 rData2[24]
port 70 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 rData2[25]
port 71 nsew signal output
rlabel metal2 s 215114 0 215170 800 6 rData2[26]
port 72 nsew signal output
rlabel metal3 s 243523 38088 244323 38208 6 rData2[27]
port 73 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 rData2[28]
port 74 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 rData2[29]
port 75 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 rData2[2]
port 76 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 rData2[30]
port 77 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 rData2[31]
port 78 nsew signal output
rlabel metal3 s 243523 168648 244323 168768 6 rData2[3]
port 79 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 rData2[4]
port 80 nsew signal output
rlabel metal2 s 235078 0 235134 800 6 rData2[5]
port 81 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 rData2[6]
port 82 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 rData2[7]
port 83 nsew signal output
rlabel metal2 s 136546 185138 136602 185938 6 rData2[8]
port 84 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 rData2[9]
port 85 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 reset
port 86 nsew signal input
rlabel metal4 s 4208 2128 4528 183376 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 183376 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 183376 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 183376 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 183376 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 183376 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 183376 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 183376 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 183376 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 183376 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 183376 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 183376 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 183376 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 183376 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 183376 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 183376 6 vssd1
port 88 nsew ground bidirectional
rlabel metal2 s 77942 0 77998 800 6 wAddr1[0]
port 89 nsew signal input
rlabel metal2 s 227994 0 228050 800 6 wAddr1[1]
port 90 nsew signal input
rlabel metal3 s 243523 113568 244323 113688 6 wAddr1[2]
port 91 nsew signal input
rlabel metal3 s 243523 65288 244323 65408 6 wAddr1[3]
port 92 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 wAddr1[4]
port 93 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 wAddr2[0]
port 94 nsew signal input
rlabel metal3 s 243523 17008 244323 17128 6 wAddr2[1]
port 95 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 wAddr2[2]
port 96 nsew signal input
rlabel metal3 s 243523 78888 244323 79008 6 wAddr2[3]
port 97 nsew signal input
rlabel metal3 s 243523 141448 244323 141568 6 wAddr2[4]
port 98 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 wData[0]
port 99 nsew signal input
rlabel metal3 s 243523 155048 244323 155168 6 wData[10]
port 100 nsew signal input
rlabel metal2 s 12898 185138 12954 185938 6 wData[11]
port 101 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 wData[12]
port 102 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 wData[13]
port 103 nsew signal input
rlabel metal2 s 18 0 74 800 6 wData[14]
port 104 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 wData[15]
port 105 nsew signal input
rlabel metal2 s 32218 185138 32274 185938 6 wData[16]
port 106 nsew signal input
rlabel metal2 s 97262 185138 97318 185938 6 wData[17]
port 107 nsew signal input
rlabel metal2 s 169390 185138 169446 185938 6 wData[18]
port 108 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 wData[19]
port 109 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 wData[1]
port 110 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wData[20]
port 111 nsew signal input
rlabel metal2 s 202234 185138 202290 185938 6 wData[21]
port 112 nsew signal input
rlabel metal2 s 156510 185138 156566 185938 6 wData[22]
port 113 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 wData[23]
port 114 nsew signal input
rlabel metal2 s 227994 185138 228050 185938 6 wData[24]
port 115 nsew signal input
rlabel metal3 s 243523 3408 244323 3528 6 wData[25]
port 116 nsew signal input
rlabel metal2 s 19338 185138 19394 185938 6 wData[26]
port 117 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 wData[27]
port 118 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wData[28]
port 119 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 wData[29]
port 120 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 wData[2]
port 121 nsew signal input
rlabel metal3 s 243523 106768 244323 106888 6 wData[30]
port 122 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 wData[31]
port 123 nsew signal input
rlabel metal2 s 195150 185138 195206 185938 6 wData[3]
port 124 nsew signal input
rlabel metal2 s 188710 185138 188766 185938 6 wData[4]
port 125 nsew signal input
rlabel metal2 s 38658 185138 38714 185938 6 wData[5]
port 126 nsew signal input
rlabel metal2 s 71502 185138 71558 185938 6 wData[6]
port 127 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 wData[7]
port 128 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 wData[8]
port 129 nsew signal input
rlabel metal2 s 5814 185138 5870 185938 6 wData[9]
port 130 nsew signal input
rlabel metal3 s 243523 72088 244323 72208 6 wEnable
port 131 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 244323 185938
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 109227966
string GDS_FILE /home/courtney/Desktop/Caravel-Vector-Coprocessor-AI/openlane/VectorRegFile/runs/23_08_17_12_46/results/signoff/VectorRegFile.magic.gds
string GDS_START 606374
<< end >>

