magic
tech sky130A
magscale 1 2
timestamp 1692640444
<< metal1 >>
rect 19058 684020 19064 684072
rect 19116 684060 19122 684072
rect 43898 684060 43904 684072
rect 19116 684032 43904 684060
rect 19116 684020 19122 684032
rect 43898 684020 43904 684032
rect 43956 684020 43962 684072
rect 19150 683952 19156 684004
rect 19208 683992 19214 684004
rect 65794 683992 65800 684004
rect 19208 683964 65800 683992
rect 19208 683952 19214 683964
rect 65794 683952 65800 683964
rect 65852 683952 65858 684004
rect 15930 683884 15936 683936
rect 15988 683924 15994 683936
rect 87046 683924 87052 683936
rect 15988 683896 87052 683924
rect 15988 683884 15994 683896
rect 87046 683884 87052 683896
rect 87104 683884 87110 683936
rect 17494 683816 17500 683868
rect 17552 683856 17558 683868
rect 108942 683856 108948 683868
rect 17552 683828 108948 683856
rect 17552 683816 17558 683828
rect 108942 683816 108948 683828
rect 109000 683816 109006 683868
rect 21818 683748 21824 683800
rect 21876 683788 21882 683800
rect 130194 683788 130200 683800
rect 21876 683760 130200 683788
rect 21876 683748 21882 683760
rect 130194 683748 130200 683760
rect 130252 683748 130258 683800
rect 18966 683680 18972 683732
rect 19024 683720 19030 683732
rect 152090 683720 152096 683732
rect 19024 683692 152096 683720
rect 19024 683680 19030 683692
rect 152090 683680 152096 683692
rect 152148 683680 152154 683732
rect 17862 683612 17868 683664
rect 17920 683652 17926 683664
rect 173342 683652 173348 683664
rect 17920 683624 173348 683652
rect 17920 683612 17926 683624
rect 173342 683612 173348 683624
rect 173400 683612 173406 683664
rect 17770 683544 17776 683596
rect 17828 683584 17834 683596
rect 195238 683584 195244 683596
rect 17828 683556 195244 683584
rect 17828 683544 17834 683556
rect 195238 683544 195244 683556
rect 195296 683544 195302 683596
rect 18874 683476 18880 683528
rect 18932 683516 18938 683528
rect 216490 683516 216496 683528
rect 18932 683488 216496 683516
rect 18932 683476 18938 683488
rect 216490 683476 216496 683488
rect 216548 683476 216554 683528
rect 17402 683408 17408 683460
rect 17460 683448 17466 683460
rect 238386 683448 238392 683460
rect 17460 683420 238392 683448
rect 17460 683408 17466 683420
rect 238386 683408 238392 683420
rect 238444 683408 238450 683460
rect 18782 683340 18788 683392
rect 18840 683380 18846 683392
rect 259638 683380 259644 683392
rect 18840 683352 259644 683380
rect 18840 683340 18846 683352
rect 259638 683340 259644 683352
rect 259696 683340 259702 683392
rect 2866 683272 2872 683324
rect 2924 683312 2930 683324
rect 302786 683312 302792 683324
rect 2924 683284 302792 683312
rect 2924 683272 2930 683284
rect 302786 683272 302792 683284
rect 302844 683272 302850 683324
rect 17586 683204 17592 683256
rect 17644 683244 17650 683256
rect 389082 683244 389088 683256
rect 17644 683216 389088 683244
rect 17644 683204 17650 683216
rect 389082 683204 389088 683216
rect 389140 683204 389146 683256
rect 540422 683204 540428 683256
rect 540480 683244 540486 683256
rect 564434 683244 564440 683256
rect 540480 683216 564440 683244
rect 540480 683204 540486 683216
rect 564434 683204 564440 683216
rect 564492 683204 564498 683256
rect 19242 683136 19248 683188
rect 19300 683176 19306 683188
rect 454126 683176 454132 683188
rect 19300 683148 454132 683176
rect 19300 683136 19306 683148
rect 454126 683136 454132 683148
rect 454184 683136 454190 683188
rect 497274 683136 497280 683188
rect 497332 683176 497338 683188
rect 564526 683176 564532 683188
rect 497332 683148 564532 683176
rect 497332 683136 497338 683148
rect 564526 683136 564532 683148
rect 564584 683136 564590 683188
rect 307754 681572 307760 681624
rect 307812 681612 307818 681624
rect 307812 681584 312860 681612
rect 307812 681572 307818 681584
rect 312538 681544 312544 681556
rect 311636 681516 312544 681544
rect 307708 681368 307714 681420
rect 307766 681368 307772 681420
rect 20530 681300 20536 681352
rect 20588 681340 20594 681352
rect 307726 681340 307754 681368
rect 20588 681312 307754 681340
rect 20588 681300 20594 681312
rect 8754 681232 8760 681284
rect 8812 681272 8818 681284
rect 311636 681272 311664 681516
rect 312538 681504 312544 681516
rect 312596 681504 312602 681556
rect 312832 681476 312860 681584
rect 8812 681244 311664 681272
rect 311728 681448 312676 681476
rect 312832 681448 325694 681476
rect 8812 681232 8818 681244
rect 566 681164 572 681216
rect 624 681204 630 681216
rect 311728 681204 311756 681448
rect 312538 681368 312544 681420
rect 312596 681368 312602 681420
rect 312648 681408 312676 681448
rect 324406 681408 324412 681420
rect 312648 681380 324412 681408
rect 324406 681368 324412 681380
rect 324464 681368 324470 681420
rect 624 681176 311756 681204
rect 312556 681204 312584 681368
rect 325666 681340 325694 681448
rect 518158 681408 518164 681420
rect 509206 681380 518164 681408
rect 509206 681340 509234 681380
rect 518158 681368 518164 681380
rect 518216 681368 518222 681420
rect 325666 681312 509234 681340
rect 561858 681272 561864 681284
rect 325666 681244 561864 681272
rect 325666 681204 325694 681244
rect 561858 681232 561864 681244
rect 561916 681232 561922 681284
rect 312556 681176 325694 681204
rect 624 681164 630 681176
rect 11146 659676 11152 659728
rect 11204 659716 11210 659728
rect 19334 659716 19340 659728
rect 11204 659688 19340 659716
rect 11204 659676 11210 659688
rect 19334 659676 19340 659688
rect 19392 659676 19398 659728
rect 18230 614116 18236 614168
rect 18288 614156 18294 614168
rect 20162 614156 20168 614168
rect 18288 614128 20168 614156
rect 18288 614116 18294 614128
rect 20162 614116 20168 614128
rect 20220 614116 20226 614168
rect 5258 545096 5264 545148
rect 5316 545136 5322 545148
rect 19334 545136 19340 545148
rect 5316 545108 19340 545136
rect 5316 545096 5322 545108
rect 19334 545096 19340 545108
rect 19392 545096 19398 545148
rect 14458 499536 14464 499588
rect 14516 499576 14522 499588
rect 19334 499576 19340 499588
rect 14516 499548 19340 499576
rect 14516 499536 14522 499548
rect 19334 499536 19340 499548
rect 19392 499536 19398 499588
rect 1670 454656 1676 454708
rect 1728 454696 1734 454708
rect 19702 454696 19708 454708
rect 1728 454668 19708 454696
rect 1728 454656 1734 454668
rect 19702 454656 19708 454668
rect 19760 454656 19766 454708
rect 7650 271872 7656 271924
rect 7708 271912 7714 271924
rect 19334 271912 19340 271924
rect 7708 271884 19340 271912
rect 7708 271872 7714 271884
rect 19334 271872 19340 271884
rect 19392 271872 19398 271924
rect 17218 135260 17224 135312
rect 17276 135300 17282 135312
rect 19518 135300 19524 135312
rect 17276 135272 19524 135300
rect 17276 135260 17282 135272
rect 19518 135260 19524 135272
rect 19576 135260 19582 135312
rect 17310 22788 17316 22840
rect 17368 22828 17374 22840
rect 17368 22800 33456 22828
rect 17368 22788 17374 22800
rect 18690 22720 18696 22772
rect 18748 22760 18754 22772
rect 18748 22732 26234 22760
rect 18748 22720 18754 22732
rect 26206 22692 26234 22732
rect 26206 22664 33364 22692
rect 33336 22488 33364 22664
rect 33428 22624 33456 22800
rect 36280 22732 38654 22760
rect 36280 22636 36308 22732
rect 38626 22692 38654 22732
rect 43180 22732 45554 22760
rect 43180 22692 43208 22732
rect 38626 22664 43208 22692
rect 33428 22596 33548 22624
rect 33520 22556 33548 22596
rect 36262 22584 36268 22636
rect 36320 22584 36326 22636
rect 43070 22624 43076 22636
rect 38626 22596 43076 22624
rect 38626 22556 38654 22596
rect 43070 22584 43076 22596
rect 43128 22584 43134 22636
rect 45526 22624 45554 22732
rect 46658 22624 46664 22636
rect 45526 22596 46664 22624
rect 46658 22584 46664 22596
rect 46716 22584 46722 22636
rect 33520 22528 38654 22556
rect 36262 22488 36268 22500
rect 33336 22460 36268 22488
rect 36262 22448 36268 22460
rect 36320 22448 36326 22500
rect 18966 21972 18972 22024
rect 19024 22012 19030 22024
rect 52546 22012 52552 22024
rect 19024 21984 52552 22012
rect 19024 21972 19030 21984
rect 52546 21972 52552 21984
rect 52604 21972 52610 22024
rect 18874 21904 18880 21956
rect 18932 21944 18938 21956
rect 58434 21944 58440 21956
rect 18932 21916 58440 21944
rect 18932 21904 18938 21916
rect 58434 21904 58440 21916
rect 58492 21904 58498 21956
rect 17862 21836 17868 21888
rect 17920 21876 17926 21888
rect 59630 21876 59636 21888
rect 17920 21848 59636 21876
rect 17920 21836 17926 21848
rect 59630 21836 59636 21848
rect 59688 21836 59694 21888
rect 18782 21768 18788 21820
rect 18840 21808 18846 21820
rect 65518 21808 65524 21820
rect 18840 21780 65524 21808
rect 18840 21768 18846 21780
rect 65518 21768 65524 21780
rect 65576 21768 65582 21820
rect 17770 21700 17776 21752
rect 17828 21740 17834 21752
rect 73798 21740 73804 21752
rect 17828 21712 73804 21740
rect 17828 21700 17834 21712
rect 73798 21700 73804 21712
rect 73856 21700 73862 21752
rect 17494 21632 17500 21684
rect 17552 21672 17558 21684
rect 84470 21672 84476 21684
rect 17552 21644 84476 21672
rect 17552 21632 17558 21644
rect 84470 21632 84476 21644
rect 84528 21632 84534 21684
rect 17586 21564 17592 21616
rect 17644 21604 17650 21616
rect 86862 21604 86868 21616
rect 17644 21576 86868 21604
rect 17644 21564 17650 21576
rect 86862 21564 86868 21576
rect 86920 21564 86926 21616
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 89162 21536 89168 21548
rect 17460 21508 89168 21536
rect 17460 21496 17466 21508
rect 89162 21496 89168 21508
rect 89220 21496 89226 21548
rect 17678 21428 17684 21480
rect 17736 21468 17742 21480
rect 90358 21468 90364 21480
rect 17736 21440 90364 21468
rect 17736 21428 17742 21440
rect 90358 21428 90364 21440
rect 90416 21428 90422 21480
rect 47854 21360 47860 21412
rect 47912 21400 47918 21412
rect 564618 21400 564624 21412
rect 47912 21372 564624 21400
rect 47912 21360 47918 21372
rect 564618 21360 564624 21372
rect 564676 21360 564682 21412
rect 28902 20612 28908 20664
rect 28960 20652 28966 20664
rect 215846 20652 215852 20664
rect 28960 20624 215852 20652
rect 28960 20612 28966 20624
rect 215846 20612 215852 20624
rect 215904 20612 215910 20664
rect 43254 20544 43260 20596
rect 43312 20584 43318 20596
rect 82170 20584 82176 20596
rect 43312 20556 82176 20584
rect 43312 20544 43318 20556
rect 82170 20544 82176 20556
rect 82228 20544 82234 20596
rect 114002 20544 114008 20596
rect 114060 20584 114066 20596
rect 302142 20584 302148 20596
rect 114060 20556 302148 20584
rect 114060 20544 114066 20556
rect 302142 20544 302148 20556
rect 302200 20544 302206 20596
rect 40678 20476 40684 20528
rect 40736 20516 40742 20528
rect 237742 20516 237748 20528
rect 40736 20488 237748 20516
rect 40736 20476 40742 20488
rect 237742 20476 237748 20488
rect 237800 20476 237806 20528
rect 78582 20408 78588 20460
rect 78640 20448 78646 20460
rect 324038 20448 324044 20460
rect 78640 20420 324044 20448
rect 78640 20408 78646 20420
rect 324038 20408 324044 20420
rect 324096 20408 324102 20460
rect 39574 20340 39580 20392
rect 39632 20380 39638 20392
rect 345290 20380 345296 20392
rect 39632 20352 345296 20380
rect 39632 20340 39638 20352
rect 345290 20340 345296 20352
rect 345348 20340 345354 20392
rect 14734 20272 14740 20324
rect 14792 20312 14798 20324
rect 388438 20312 388444 20324
rect 14792 20284 388444 20312
rect 14792 20272 14798 20284
rect 388438 20272 388444 20284
rect 388496 20272 388502 20324
rect 13538 20204 13544 20256
rect 13596 20244 13602 20256
rect 65150 20244 65156 20256
rect 13596 20216 65156 20244
rect 13596 20204 13602 20216
rect 65150 20204 65156 20216
rect 65208 20204 65214 20256
rect 98638 20204 98644 20256
rect 98696 20244 98702 20256
rect 474734 20244 474740 20256
rect 98696 20216 474740 20244
rect 98696 20204 98702 20216
rect 474734 20204 474740 20216
rect 474792 20204 474798 20256
rect 23014 20136 23020 20188
rect 23072 20176 23078 20188
rect 410334 20176 410340 20188
rect 23072 20148 410340 20176
rect 23072 20136 23078 20148
rect 410334 20136 410340 20148
rect 410392 20136 410398 20188
rect 45462 20068 45468 20120
rect 45520 20108 45526 20120
rect 453482 20108 453488 20120
rect 45520 20080 453488 20108
rect 45520 20068 45526 20080
rect 453482 20068 453488 20080
rect 453540 20068 453546 20120
rect 21082 20000 21088 20052
rect 21140 20040 21146 20052
rect 431586 20040 431592 20052
rect 21140 20012 431592 20040
rect 21140 20000 21146 20012
rect 431586 20000 431592 20012
rect 431644 20000 431650 20052
rect 64322 19932 64328 19984
rect 64380 19972 64386 19984
rect 517882 19972 517888 19984
rect 64380 19944 517888 19972
rect 64380 19932 64386 19944
rect 517882 19932 517888 19944
rect 517940 19932 517946 19984
rect 102226 19864 102232 19916
rect 102284 19904 102290 19916
rect 258994 19904 259000 19916
rect 102284 19876 259000 19904
rect 102284 19864 102290 19876
rect 258994 19864 259000 19876
rect 259052 19864 259058 19916
rect 24210 19796 24216 19848
rect 24268 19836 24274 19848
rect 129550 19836 129556 19848
rect 24268 19808 129556 19836
rect 24268 19796 24274 19808
rect 129550 19796 129556 19808
rect 129608 19796 129614 19848
rect 70302 19728 70308 19780
rect 70360 19768 70366 19780
rect 172698 19768 172704 19780
rect 70360 19740 172704 19768
rect 70360 19728 70366 19740
rect 172698 19728 172704 19740
rect 172756 19728 172762 19780
rect 107010 19320 107016 19372
rect 107068 19360 107074 19372
rect 108298 19360 108304 19372
rect 107068 19332 108304 19360
rect 107068 19320 107074 19332
rect 108298 19320 108304 19332
rect 108356 19320 108362 19372
rect 76190 6808 76196 6860
rect 76248 6848 76254 6860
rect 150434 6848 150440 6860
rect 76248 6820 150440 6848
rect 76248 6808 76254 6820
rect 150434 6808 150440 6820
rect 150492 6808 150498 6860
rect 93946 6740 93952 6792
rect 94004 6780 94010 6792
rect 194594 6780 194600 6792
rect 94004 6752 194600 6780
rect 94004 6740 94010 6752
rect 194594 6740 194600 6752
rect 194652 6740 194658 6792
rect 115198 6672 115204 6724
rect 115256 6712 115262 6724
rect 367094 6712 367100 6724
rect 115256 6684 367100 6712
rect 115256 6672 115262 6684
rect 367094 6672 367100 6684
rect 367152 6672 367158 6724
rect 116394 6604 116400 6656
rect 116452 6644 116458 6656
rect 562502 6644 562508 6656
rect 116452 6616 562508 6644
rect 116452 6604 116458 6616
rect 562502 6604 562508 6616
rect 562560 6604 562566 6656
rect 87966 6536 87972 6588
rect 88024 6576 88030 6588
rect 562410 6576 562416 6588
rect 88024 6548 562416 6576
rect 88024 6536 88030 6548
rect 562410 6536 562416 6548
rect 562468 6536 562474 6588
rect 19794 6468 19800 6520
rect 19852 6508 19858 6520
rect 66714 6508 66720 6520
rect 19852 6480 66720 6508
rect 19852 6468 19858 6480
rect 66714 6468 66720 6480
rect 66772 6468 66778 6520
rect 77386 6468 77392 6520
rect 77444 6508 77450 6520
rect 563882 6508 563888 6520
rect 77444 6480 563888 6508
rect 77444 6468 77450 6480
rect 563882 6468 563888 6480
rect 563940 6468 563946 6520
rect 63218 6400 63224 6452
rect 63276 6440 63282 6452
rect 561858 6440 561864 6452
rect 63276 6412 561864 6440
rect 63276 6400 63282 6412
rect 561858 6400 561864 6412
rect 561916 6400 561922 6452
rect 56042 6332 56048 6384
rect 56100 6372 56106 6384
rect 562134 6372 562140 6384
rect 56100 6344 562140 6372
rect 56100 6332 56106 6344
rect 562134 6332 562140 6344
rect 562192 6332 562198 6384
rect 38378 6264 38384 6316
rect 38436 6304 38442 6316
rect 562042 6304 562048 6316
rect 38436 6276 562048 6304
rect 38436 6264 38442 6276
rect 562042 6264 562048 6276
rect 562100 6264 562106 6316
rect 34790 6196 34796 6248
rect 34848 6236 34854 6248
rect 562594 6236 562600 6248
rect 34848 6208 562600 6236
rect 34848 6196 34854 6208
rect 562594 6196 562600 6208
rect 562652 6196 562658 6248
rect 12342 6128 12348 6180
rect 12400 6168 12406 6180
rect 560294 6168 560300 6180
rect 12400 6140 560300 6168
rect 12400 6128 12406 6140
rect 560294 6128 560300 6140
rect 560352 6128 560358 6180
rect 21266 5380 21272 5432
rect 21324 5420 21330 5432
rect 44266 5420 44272 5432
rect 21324 5392 44272 5420
rect 21324 5380 21330 5392
rect 44266 5380 44272 5392
rect 44324 5380 44330 5432
rect 20346 5312 20352 5364
rect 20404 5352 20410 5364
rect 112806 5352 112812 5364
rect 20404 5324 112812 5352
rect 20404 5312 20410 5324
rect 112806 5312 112812 5324
rect 112864 5312 112870 5364
rect 20162 5244 20168 5296
rect 20220 5284 20226 5296
rect 108114 5284 108120 5296
rect 20220 5256 108120 5284
rect 20220 5244 20226 5256
rect 108114 5244 108120 5256
rect 108172 5244 108178 5296
rect 111610 5244 111616 5296
rect 111668 5284 111674 5296
rect 280154 5284 280160 5296
rect 111668 5256 280160 5284
rect 111668 5244 111674 5256
rect 280154 5244 280160 5256
rect 280212 5244 280218 5296
rect 20530 5176 20536 5228
rect 20588 5216 20594 5228
rect 83274 5216 83280 5228
rect 20588 5188 83280 5216
rect 20588 5176 20594 5188
rect 83274 5176 83280 5188
rect 83332 5176 83338 5228
rect 97442 5176 97448 5228
rect 97500 5216 97506 5228
rect 539594 5216 539600 5228
rect 97500 5188 539600 5216
rect 97500 5176 97506 5188
rect 539594 5176 539600 5188
rect 539652 5176 539658 5228
rect 19886 5108 19892 5160
rect 19944 5148 19950 5160
rect 118602 5148 118608 5160
rect 19944 5120 118608 5148
rect 19944 5108 19950 5120
rect 118602 5108 118608 5120
rect 118660 5108 118666 5160
rect 118694 5108 118700 5160
rect 118752 5148 118758 5160
rect 563514 5148 563520 5160
rect 118752 5120 563520 5148
rect 118752 5108 118758 5120
rect 563514 5108 563520 5120
rect 563572 5108 563578 5160
rect 19978 5040 19984 5092
rect 20036 5080 20042 5092
rect 92750 5080 92756 5092
rect 20036 5052 92756 5080
rect 20036 5040 20042 5052
rect 92750 5040 92756 5052
rect 92808 5040 92814 5092
rect 104526 5040 104532 5092
rect 104584 5080 104590 5092
rect 562318 5080 562324 5092
rect 104584 5052 562324 5080
rect 104584 5040 104590 5052
rect 562318 5040 562324 5052
rect 562376 5040 562382 5092
rect 21174 4972 21180 5024
rect 21232 5012 21238 5024
rect 48958 5012 48964 5024
rect 21232 4984 48964 5012
rect 21232 4972 21238 4984
rect 48958 4972 48964 4984
rect 49016 4972 49022 5024
rect 80882 4972 80888 5024
rect 80940 5012 80946 5024
rect 561950 5012 561956 5024
rect 80940 4984 561956 5012
rect 80940 4972 80946 4984
rect 561950 4972 561956 4984
rect 562008 4972 562014 5024
rect 20438 4904 20444 4956
rect 20496 4944 20502 4956
rect 69106 4944 69112 4956
rect 20496 4916 69112 4944
rect 20496 4904 20502 4916
rect 69106 4904 69112 4916
rect 69164 4904 69170 4956
rect 72602 4904 72608 4956
rect 72660 4944 72666 4956
rect 562226 4944 562232 4956
rect 72660 4916 562232 4944
rect 72660 4904 72666 4916
rect 562226 4904 562232 4916
rect 562284 4904 562290 4956
rect 21818 4836 21824 4888
rect 21876 4876 21882 4888
rect 563698 4876 563704 4888
rect 21876 4848 563704 4876
rect 21876 4836 21882 4848
rect 563698 4836 563704 4848
rect 563756 4836 563762 4888
rect 17034 4768 17040 4820
rect 17092 4808 17098 4820
rect 563606 4808 563612 4820
rect 17092 4780 563612 4808
rect 17092 4768 17098 4780
rect 563606 4768 563612 4780
rect 563664 4768 563670 4820
rect 18598 4088 18604 4140
rect 18656 4128 18662 4140
rect 62022 4128 62028 4140
rect 18656 4100 62028 4128
rect 18656 4088 18662 4100
rect 62022 4088 62028 4100
rect 62080 4088 62086 4140
rect 21910 4020 21916 4072
rect 21968 4060 21974 4072
rect 71498 4060 71504 4072
rect 21968 4032 71504 4060
rect 21968 4020 21974 4032
rect 71498 4020 71504 4032
rect 71556 4020 71562 4072
rect 19058 3952 19064 4004
rect 19116 3992 19122 4004
rect 74994 3992 75000 4004
rect 19116 3964 75000 3992
rect 19116 3952 19122 3964
rect 74994 3952 75000 3964
rect 75052 3952 75058 4004
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 85574 3924 85580 3936
rect 27764 3896 85580 3924
rect 27764 3884 27770 3896
rect 85574 3884 85580 3896
rect 85632 3884 85638 3936
rect 119890 3884 119896 3936
rect 119948 3924 119954 3936
rect 495434 3924 495440 3936
rect 119948 3896 495440 3924
rect 119948 3884 119954 3896
rect 495434 3884 495440 3896
rect 495492 3884 495498 3936
rect 22002 3816 22008 3868
rect 22060 3856 22066 3868
rect 82078 3856 82084 3868
rect 22060 3828 82084 3856
rect 22060 3816 22066 3828
rect 82078 3816 82084 3828
rect 82136 3816 82142 3868
rect 82170 3816 82176 3868
rect 82228 3856 82234 3868
rect 103330 3856 103336 3868
rect 82228 3828 103336 3856
rect 82228 3816 82234 3828
rect 103330 3816 103336 3828
rect 103388 3816 103394 3868
rect 105722 3816 105728 3868
rect 105780 3856 105786 3868
rect 118694 3856 118700 3868
rect 105780 3828 118700 3856
rect 105780 3816 105786 3828
rect 118694 3816 118700 3828
rect 118752 3816 118758 3868
rect 124674 3816 124680 3868
rect 124732 3856 124738 3868
rect 563146 3856 563152 3868
rect 124732 3828 563152 3856
rect 124732 3816 124738 3828
rect 563146 3816 563152 3828
rect 563204 3816 563210 3868
rect 19150 3748 19156 3800
rect 19208 3788 19214 3800
rect 85666 3788 85672 3800
rect 19208 3760 85672 3788
rect 19208 3748 19214 3760
rect 85666 3748 85672 3760
rect 85724 3748 85730 3800
rect 99834 3748 99840 3800
rect 99892 3788 99898 3800
rect 107010 3788 107016 3800
rect 99892 3760 107016 3788
rect 99892 3748 99898 3760
rect 107010 3748 107016 3760
rect 107068 3748 107074 3800
rect 117590 3748 117596 3800
rect 117648 3788 117654 3800
rect 564434 3788 564440 3800
rect 117648 3760 564440 3788
rect 117648 3748 117654 3760
rect 564434 3748 564440 3760
rect 564492 3748 564498 3800
rect 21358 3680 21364 3732
rect 21416 3720 21422 3732
rect 21416 3692 21496 3720
rect 21416 3680 21422 3692
rect 17218 3612 17224 3664
rect 17276 3652 17282 3664
rect 21468 3652 21496 3692
rect 21634 3680 21640 3732
rect 21692 3720 21698 3732
rect 96246 3720 96252 3732
rect 21692 3692 96252 3720
rect 21692 3680 21698 3692
rect 96246 3680 96252 3692
rect 96304 3680 96310 3732
rect 106918 3680 106924 3732
rect 106976 3720 106982 3732
rect 564526 3720 564532 3732
rect 106976 3692 564532 3720
rect 106976 3680 106982 3692
rect 564526 3680 564532 3692
rect 564584 3680 564590 3732
rect 53742 3652 53748 3664
rect 17276 3624 21404 3652
rect 21468 3624 53748 3652
rect 17276 3612 17282 3624
rect 20254 3544 20260 3596
rect 20312 3584 20318 3596
rect 21376 3584 21404 3624
rect 53742 3612 53748 3624
rect 53800 3612 53806 3664
rect 60826 3612 60832 3664
rect 60884 3652 60890 3664
rect 563054 3652 563060 3664
rect 60884 3624 563060 3652
rect 60884 3612 60890 3624
rect 563054 3612 563060 3624
rect 563112 3612 563118 3664
rect 51350 3584 51356 3596
rect 20312 3556 21312 3584
rect 21376 3556 51356 3584
rect 20312 3544 20318 3556
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 14458 3516 14464 3528
rect 10008 3488 14464 3516
rect 10008 3476 10014 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 21082 3516 21088 3528
rect 20680 3488 21088 3516
rect 20680 3476 20686 3488
rect 21082 3476 21088 3488
rect 21140 3476 21146 3528
rect 21284 3516 21312 3556
rect 51350 3544 51356 3556
rect 51408 3544 51414 3596
rect 57238 3544 57244 3596
rect 57296 3584 57302 3596
rect 563330 3584 563336 3596
rect 57296 3556 563336 3584
rect 57296 3544 57302 3556
rect 563330 3544 563336 3556
rect 563388 3544 563394 3596
rect 31294 3516 31300 3528
rect 21284 3488 31300 3516
rect 31294 3476 31300 3488
rect 31352 3476 31358 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 563422 3516 563428 3528
rect 41932 3488 563428 3516
rect 41932 3476 41938 3488
rect 563422 3476 563428 3488
rect 563480 3476 563486 3528
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 563790 3448 563796 3460
rect 19484 3420 563796 3448
rect 19484 3408 19490 3420
rect 563790 3408 563796 3420
rect 563848 3408 563854 3460
rect 21542 3340 21548 3392
rect 21600 3380 21606 3392
rect 50154 3380 50160 3392
rect 21600 3352 50160 3380
rect 21600 3340 21606 3352
rect 50154 3340 50160 3352
rect 50212 3340 50218 3392
rect 21450 3272 21456 3324
rect 21508 3312 21514 3324
rect 32398 3312 32404 3324
rect 21508 3284 32404 3312
rect 21508 3272 21514 3284
rect 32398 3272 32404 3284
rect 32456 3272 32462 3324
rect 20530 3204 20536 3256
rect 20588 3244 20594 3256
rect 30098 3244 30104 3256
rect 20588 3216 30104 3244
rect 20588 3204 20594 3216
rect 30098 3204 30104 3216
rect 30156 3204 30162 3256
rect 20070 2864 20076 2916
rect 20128 2904 20134 2916
rect 25314 2904 25320 2916
rect 20128 2876 25320 2904
rect 20128 2864 20134 2876
rect 25314 2864 25320 2876
rect 25372 2864 25378 2916
<< via1 >>
rect 19064 684020 19116 684072
rect 43904 684020 43956 684072
rect 19156 683952 19208 684004
rect 65800 683952 65852 684004
rect 15936 683884 15988 683936
rect 87052 683884 87104 683936
rect 17500 683816 17552 683868
rect 108948 683816 109000 683868
rect 21824 683748 21876 683800
rect 130200 683748 130252 683800
rect 18972 683680 19024 683732
rect 152096 683680 152148 683732
rect 17868 683612 17920 683664
rect 173348 683612 173400 683664
rect 17776 683544 17828 683596
rect 195244 683544 195296 683596
rect 18880 683476 18932 683528
rect 216496 683476 216548 683528
rect 17408 683408 17460 683460
rect 238392 683408 238444 683460
rect 18788 683340 18840 683392
rect 259644 683340 259696 683392
rect 2872 683272 2924 683324
rect 302792 683272 302844 683324
rect 17592 683204 17644 683256
rect 389088 683204 389140 683256
rect 540428 683204 540480 683256
rect 564440 683204 564492 683256
rect 19248 683136 19300 683188
rect 454132 683136 454184 683188
rect 497280 683136 497332 683188
rect 564532 683136 564584 683188
rect 307760 681572 307812 681624
rect 307714 681368 307766 681420
rect 20536 681300 20588 681352
rect 8760 681232 8812 681284
rect 312544 681504 312596 681556
rect 572 681164 624 681216
rect 312544 681368 312596 681420
rect 324412 681368 324464 681420
rect 518164 681368 518216 681420
rect 561864 681232 561916 681284
rect 11152 659676 11204 659728
rect 19340 659676 19392 659728
rect 18236 614116 18288 614168
rect 20168 614116 20220 614168
rect 5264 545096 5316 545148
rect 19340 545096 19392 545148
rect 14464 499536 14516 499588
rect 19340 499536 19392 499588
rect 1676 454656 1728 454708
rect 19708 454656 19760 454708
rect 7656 271872 7708 271924
rect 19340 271872 19392 271924
rect 17224 135260 17276 135312
rect 19524 135260 19576 135312
rect 17316 22788 17368 22840
rect 18696 22720 18748 22772
rect 36268 22584 36320 22636
rect 43076 22584 43128 22636
rect 46664 22584 46716 22636
rect 36268 22448 36320 22500
rect 18972 21972 19024 22024
rect 52552 21972 52604 22024
rect 18880 21904 18932 21956
rect 58440 21904 58492 21956
rect 17868 21836 17920 21888
rect 59636 21836 59688 21888
rect 18788 21768 18840 21820
rect 65524 21768 65576 21820
rect 17776 21700 17828 21752
rect 73804 21700 73856 21752
rect 17500 21632 17552 21684
rect 84476 21632 84528 21684
rect 17592 21564 17644 21616
rect 86868 21564 86920 21616
rect 17408 21496 17460 21548
rect 89168 21496 89220 21548
rect 17684 21428 17736 21480
rect 90364 21428 90416 21480
rect 47860 21360 47912 21412
rect 564624 21360 564676 21412
rect 28908 20612 28960 20664
rect 215852 20612 215904 20664
rect 43260 20544 43312 20596
rect 82176 20544 82228 20596
rect 114008 20544 114060 20596
rect 302148 20544 302200 20596
rect 40684 20476 40736 20528
rect 237748 20476 237800 20528
rect 78588 20408 78640 20460
rect 324044 20408 324096 20460
rect 39580 20340 39632 20392
rect 345296 20340 345348 20392
rect 14740 20272 14792 20324
rect 388444 20272 388496 20324
rect 13544 20204 13596 20256
rect 65156 20204 65208 20256
rect 98644 20204 98696 20256
rect 474740 20204 474792 20256
rect 23020 20136 23072 20188
rect 410340 20136 410392 20188
rect 45468 20068 45520 20120
rect 453488 20068 453540 20120
rect 21088 20000 21140 20052
rect 431592 20000 431644 20052
rect 64328 19932 64380 19984
rect 517888 19932 517940 19984
rect 102232 19864 102284 19916
rect 259000 19864 259052 19916
rect 24216 19796 24268 19848
rect 129556 19796 129608 19848
rect 70308 19728 70360 19780
rect 172704 19728 172756 19780
rect 107016 19320 107068 19372
rect 108304 19320 108356 19372
rect 76196 6808 76248 6860
rect 150440 6808 150492 6860
rect 93952 6740 94004 6792
rect 194600 6740 194652 6792
rect 115204 6672 115256 6724
rect 367100 6672 367152 6724
rect 116400 6604 116452 6656
rect 562508 6604 562560 6656
rect 87972 6536 88024 6588
rect 562416 6536 562468 6588
rect 19800 6468 19852 6520
rect 66720 6468 66772 6520
rect 77392 6468 77444 6520
rect 563888 6468 563940 6520
rect 63224 6400 63276 6452
rect 561864 6400 561916 6452
rect 56048 6332 56100 6384
rect 562140 6332 562192 6384
rect 38384 6264 38436 6316
rect 562048 6264 562100 6316
rect 34796 6196 34848 6248
rect 562600 6196 562652 6248
rect 12348 6128 12400 6180
rect 560300 6128 560352 6180
rect 21272 5380 21324 5432
rect 44272 5380 44324 5432
rect 20352 5312 20404 5364
rect 112812 5312 112864 5364
rect 20168 5244 20220 5296
rect 108120 5244 108172 5296
rect 111616 5244 111668 5296
rect 280160 5244 280212 5296
rect 20536 5176 20588 5228
rect 83280 5176 83332 5228
rect 97448 5176 97500 5228
rect 539600 5176 539652 5228
rect 19892 5108 19944 5160
rect 118608 5108 118660 5160
rect 118700 5108 118752 5160
rect 563520 5108 563572 5160
rect 19984 5040 20036 5092
rect 92756 5040 92808 5092
rect 104532 5040 104584 5092
rect 562324 5040 562376 5092
rect 21180 4972 21232 5024
rect 48964 4972 49016 5024
rect 80888 4972 80940 5024
rect 561956 4972 562008 5024
rect 20444 4904 20496 4956
rect 69112 4904 69164 4956
rect 72608 4904 72660 4956
rect 562232 4904 562284 4956
rect 21824 4836 21876 4888
rect 563704 4836 563756 4888
rect 17040 4768 17092 4820
rect 563612 4768 563664 4820
rect 18604 4088 18656 4140
rect 62028 4088 62080 4140
rect 21916 4020 21968 4072
rect 71504 4020 71556 4072
rect 19064 3952 19116 4004
rect 75000 3952 75052 4004
rect 27712 3884 27764 3936
rect 85580 3884 85632 3936
rect 119896 3884 119948 3936
rect 495440 3884 495492 3936
rect 22008 3816 22060 3868
rect 82084 3816 82136 3868
rect 82176 3816 82228 3868
rect 103336 3816 103388 3868
rect 105728 3816 105780 3868
rect 118700 3816 118752 3868
rect 124680 3816 124732 3868
rect 563152 3816 563204 3868
rect 19156 3748 19208 3800
rect 85672 3748 85724 3800
rect 99840 3748 99892 3800
rect 107016 3748 107068 3800
rect 117596 3748 117648 3800
rect 564440 3748 564492 3800
rect 21364 3680 21416 3732
rect 17224 3612 17276 3664
rect 21640 3680 21692 3732
rect 96252 3680 96304 3732
rect 106924 3680 106976 3732
rect 564532 3680 564584 3732
rect 20260 3544 20312 3596
rect 53748 3612 53800 3664
rect 60832 3612 60884 3664
rect 563060 3612 563112 3664
rect 9956 3476 10008 3528
rect 14464 3476 14516 3528
rect 20628 3476 20680 3528
rect 21088 3476 21140 3528
rect 51356 3544 51408 3596
rect 57244 3544 57296 3596
rect 563336 3544 563388 3596
rect 31300 3476 31352 3528
rect 41880 3476 41932 3528
rect 563428 3476 563480 3528
rect 19432 3408 19484 3460
rect 563796 3408 563848 3460
rect 21548 3340 21600 3392
rect 50160 3340 50212 3392
rect 21456 3272 21508 3324
rect 32404 3272 32456 3324
rect 20536 3204 20588 3256
rect 30104 3204 30156 3256
rect 20076 2864 20128 2916
rect 25320 2864 25372 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 19064 684072 19116 684078
rect 19064 684014 19116 684020
rect 43904 684072 43956 684078
rect 43904 684014 43956 684020
rect 15936 683936 15988 683942
rect 15936 683878 15988 683884
rect 2872 683324 2924 683330
rect 2872 683266 2924 683272
rect 572 681216 624 681222
rect 572 681158 624 681164
rect 584 480 612 681158
rect 1676 454708 1728 454714
rect 1676 454650 1728 454656
rect 1688 480 1716 454650
rect 2884 480 2912 683266
rect 8760 681284 8812 681290
rect 8760 681226 8812 681232
rect 5264 545148 5316 545154
rect 5264 545090 5316 545096
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4080 480 4108 6151
rect 5276 480 5304 545090
rect 7656 271924 7708 271930
rect 7656 271866 7708 271872
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 271866
rect 8772 480 8800 681226
rect 11152 659728 11204 659734
rect 11152 659670 11204 659676
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9968 480 9996 3470
rect 11164 480 11192 659670
rect 14464 499588 14516 499594
rect 14464 499530 14516 499536
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12360 480 12388 6122
rect 13556 480 13584 20198
rect 14476 3534 14504 499530
rect 14740 20324 14792 20330
rect 14740 20266 14792 20272
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14752 480 14780 20266
rect 15948 480 15976 683878
rect 17500 683868 17552 683874
rect 17500 683810 17552 683816
rect 17314 683496 17370 683505
rect 17314 683431 17370 683440
rect 17408 683460 17460 683466
rect 17224 135312 17276 135318
rect 17224 135254 17276 135260
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17052 480 17080 4762
rect 17236 3670 17264 135254
rect 17328 22846 17356 683431
rect 17408 683402 17460 683408
rect 17316 22840 17368 22846
rect 17316 22782 17368 22788
rect 17420 21554 17448 683402
rect 17512 21690 17540 683810
rect 18972 683732 19024 683738
rect 18972 683674 19024 683680
rect 17868 683664 17920 683670
rect 17868 683606 17920 683612
rect 18694 683632 18750 683641
rect 17776 683596 17828 683602
rect 17776 683538 17828 683544
rect 17682 683360 17738 683369
rect 17682 683295 17738 683304
rect 17592 683256 17644 683262
rect 17592 683198 17644 683204
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17604 21622 17632 683198
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17696 21486 17724 683295
rect 17788 21758 17816 683538
rect 17880 21894 17908 683606
rect 18694 683567 18750 683576
rect 18236 614168 18288 614174
rect 18236 614110 18288 614116
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17776 21752 17828 21758
rect 17776 21694 17828 21700
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 18248 480 18276 614110
rect 18602 363488 18658 363497
rect 18602 363423 18658 363432
rect 18616 4146 18644 363423
rect 18708 22778 18736 683567
rect 18880 683528 18932 683534
rect 18880 683470 18932 683476
rect 18788 683392 18840 683398
rect 18788 683334 18840 683340
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18800 21826 18828 683334
rect 18892 21962 18920 683470
rect 18984 22030 19012 683674
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18788 21820 18840 21826
rect 18788 21762 18840 21768
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 19076 4010 19104 684014
rect 19156 684004 19208 684010
rect 19156 683946 19208 683952
rect 19064 4004 19116 4010
rect 19064 3946 19116 3952
rect 19168 3806 19196 683946
rect 21824 683800 21876 683806
rect 21824 683742 21876 683748
rect 19248 683188 19300 683194
rect 19248 683130 19300 683136
rect 19156 3800 19208 3806
rect 19156 3742 19208 3748
rect 19260 3233 19288 683130
rect 20536 681352 20588 681358
rect 20536 681294 20588 681300
rect 19338 659968 19394 659977
rect 19338 659903 19394 659912
rect 19352 659734 19380 659903
rect 19340 659728 19392 659734
rect 19340 659670 19392 659676
rect 20166 614408 20222 614417
rect 20166 614343 20222 614352
rect 20180 614174 20208 614343
rect 20168 614168 20220 614174
rect 20168 614110 20220 614116
rect 19338 545728 19394 545737
rect 19338 545663 19394 545672
rect 19352 545154 19380 545663
rect 19340 545148 19392 545154
rect 19340 545090 19392 545096
rect 19338 500168 19394 500177
rect 19338 500103 19394 500112
rect 19352 499594 19380 500103
rect 19340 499588 19392 499594
rect 19340 499530 19392 499536
rect 19708 454708 19760 454714
rect 19708 454650 19760 454656
rect 19720 454617 19748 454650
rect 20548 454617 20576 681294
rect 21730 636848 21786 636857
rect 21730 636783 21786 636792
rect 21638 591288 21694 591297
rect 21638 591223 21694 591232
rect 20626 477728 20682 477737
rect 20626 477663 20682 477672
rect 19706 454608 19762 454617
rect 19706 454543 19762 454552
rect 20534 454608 20590 454617
rect 20534 454543 20590 454552
rect 20534 409048 20590 409057
rect 20534 408983 20590 408992
rect 20442 341048 20498 341057
rect 20442 340983 20498 340992
rect 20350 317928 20406 317937
rect 20350 317863 20406 317872
rect 20258 295488 20314 295497
rect 20258 295423 20314 295432
rect 19338 272368 19394 272377
rect 19338 272303 19394 272312
rect 19352 271930 19380 272303
rect 19340 271924 19392 271930
rect 19340 271866 19392 271872
rect 20166 249928 20222 249937
rect 20166 249863 20222 249872
rect 20074 204368 20130 204377
rect 20074 204303 20130 204312
rect 19982 181248 20038 181257
rect 19982 181183 20038 181192
rect 19522 135688 19578 135697
rect 19522 135623 19578 135632
rect 19536 135318 19564 135623
rect 19524 135312 19576 135318
rect 19524 135254 19576 135260
rect 19890 113248 19946 113257
rect 19890 113183 19946 113192
rect 19798 67688 19854 67697
rect 19798 67623 19854 67632
rect 19812 6526 19840 67623
rect 19800 6520 19852 6526
rect 19800 6462 19852 6468
rect 19904 5166 19932 113183
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 19996 5098 20024 181183
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19246 3224 19302 3233
rect 19246 3159 19302 3168
rect 19444 480 19472 3402
rect 20088 2922 20116 204303
rect 20180 5302 20208 249863
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 20272 3602 20300 295423
rect 20364 5370 20392 317863
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 20456 4962 20484 340983
rect 20548 5234 20576 408983
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20640 5114 20668 477663
rect 21546 386608 21602 386617
rect 21546 386543 21602 386552
rect 21454 226808 21510 226817
rect 21454 226743 21510 226752
rect 21362 158808 21418 158817
rect 21362 158743 21418 158752
rect 21270 90128 21326 90137
rect 21270 90063 21326 90072
rect 21178 44568 21234 44577
rect 21178 44503 21234 44512
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20548 5086 20668 5114
rect 20444 4956 20496 4962
rect 20444 4898 20496 4904
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20548 3262 20576 5086
rect 21100 3534 21128 19994
rect 21192 5030 21220 44503
rect 21284 5438 21312 90063
rect 21272 5432 21324 5438
rect 21272 5374 21324 5380
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21376 3738 21404 158743
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20536 3256 20588 3262
rect 20536 3198 20588 3204
rect 20076 2916 20128 2922
rect 20076 2858 20128 2864
rect 20640 480 20668 3470
rect 21468 3330 21496 226743
rect 21560 3398 21588 386543
rect 21652 3738 21680 591223
rect 21744 3913 21772 636783
rect 21836 23497 21864 683742
rect 43916 681972 43944 684014
rect 65800 684004 65852 684010
rect 65800 683946 65852 683952
rect 65812 681972 65840 683946
rect 87052 683936 87104 683942
rect 87052 683878 87104 683884
rect 345938 683904 345994 683913
rect 87064 681972 87092 683878
rect 108948 683868 109000 683874
rect 345938 683839 345994 683848
rect 108948 683810 109000 683816
rect 108960 681972 108988 683810
rect 130200 683800 130252 683806
rect 130200 683742 130252 683748
rect 281538 683768 281594 683777
rect 130212 681972 130240 683742
rect 152096 683732 152148 683738
rect 281538 683703 281594 683712
rect 152096 683674 152148 683680
rect 152108 681972 152136 683674
rect 173348 683664 173400 683670
rect 173348 683606 173400 683612
rect 173360 681972 173388 683606
rect 195244 683596 195296 683602
rect 195244 683538 195296 683544
rect 195256 681972 195284 683538
rect 216496 683528 216548 683534
rect 216496 683470 216548 683476
rect 216508 681972 216536 683470
rect 238392 683460 238444 683466
rect 238392 683402 238444 683408
rect 238404 681972 238432 683402
rect 259644 683392 259696 683398
rect 259644 683334 259696 683340
rect 259656 681972 259684 683334
rect 281552 681972 281580 683703
rect 302792 683324 302844 683330
rect 302792 683266 302844 683272
rect 302804 681972 302832 683266
rect 324778 683224 324834 683233
rect 324778 683159 324834 683168
rect 307760 681624 307812 681630
rect 307760 681566 307812 681572
rect 307772 681442 307800 681566
rect 312544 681556 312596 681562
rect 312544 681498 312596 681504
rect 21928 681414 22678 681442
rect 307726 681426 307800 681442
rect 312556 681426 312584 681498
rect 324792 681442 324820 683159
rect 345952 681972 345980 683839
rect 410982 683632 411038 683641
rect 410982 683567 411038 683576
rect 389088 683256 389140 683262
rect 389088 683198 389140 683204
rect 389100 681972 389128 683198
rect 410996 681972 411024 683567
rect 432234 683496 432290 683505
rect 432234 683431 432290 683440
rect 432248 681972 432276 683431
rect 475382 683360 475438 683369
rect 475382 683295 475438 683304
rect 454132 683188 454184 683194
rect 454132 683130 454184 683136
rect 454144 681972 454172 683130
rect 475396 681972 475424 683295
rect 540428 683256 540480 683262
rect 540428 683198 540480 683204
rect 564440 683256 564492 683262
rect 564440 683198 564492 683204
rect 497280 683188 497332 683194
rect 497280 683130 497332 683136
rect 497292 681972 497320 683130
rect 540440 681972 540468 683198
rect 324424 681426 324820 681442
rect 518176 681426 518558 681442
rect 307714 681420 307800 681426
rect 21822 23488 21878 23497
rect 21822 23423 21878 23432
rect 21824 4888 21876 4894
rect 21824 4830 21876 4836
rect 21730 3904 21786 3913
rect 21730 3839 21786 3848
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21456 3324 21508 3330
rect 21456 3266 21508 3272
rect 21836 480 21864 4830
rect 21928 4078 21956 681414
rect 307766 681414 307800 681420
rect 312544 681420 312596 681426
rect 307714 681362 307766 681368
rect 312544 681362 312596 681368
rect 324412 681420 324820 681426
rect 324464 681414 324820 681420
rect 518164 681420 518558 681426
rect 324412 681362 324464 681368
rect 518216 681414 518558 681420
rect 518164 681362 518216 681368
rect 367834 681320 367890 681329
rect 561706 681290 561904 681306
rect 561706 681284 561916 681290
rect 561706 681278 561864 681284
rect 367834 681255 367890 681264
rect 561864 681226 561916 681232
rect 563058 679960 563114 679969
rect 563058 679895 563114 679904
rect 561862 567624 561918 567633
rect 561862 567559 561918 567568
rect 26514 22672 26570 22681
rect 26514 22607 26570 22616
rect 33598 22672 33654 22681
rect 33598 22607 33654 22616
rect 36268 22636 36320 22642
rect 21916 4072 21968 4078
rect 21916 4014 21968 4020
rect 22020 3874 22048 22100
rect 23020 20188 23072 20194
rect 23020 20130 23072 20136
rect 22008 3868 22060 3874
rect 22008 3810 22060 3816
rect 23032 480 23060 20130
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24228 480 24256 19790
rect 25320 2916 25372 2922
rect 25320 2858 25372 2864
rect 25332 480 25360 2858
rect 26528 480 26556 22607
rect 28908 20664 28960 20670
rect 28908 20606 28960 20612
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 27724 480 27752 3878
rect 28920 480 28948 20606
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 30104 3256 30156 3262
rect 30104 3198 30156 3204
rect 30116 480 30144 3198
rect 31312 480 31340 3470
rect 32404 3324 32456 3330
rect 32404 3266 32456 3272
rect 32416 480 32444 3266
rect 33612 480 33640 22607
rect 36268 22578 36320 22584
rect 43076 22636 43128 22642
rect 43076 22578 43128 22584
rect 46664 22636 46716 22642
rect 46664 22578 46716 22584
rect 36280 22506 36308 22578
rect 36268 22500 36320 22506
rect 36268 22442 36320 22448
rect 40684 20528 40736 20534
rect 40684 20470 40736 20476
rect 39580 20392 39632 20398
rect 39580 20334 39632 20340
rect 37186 6352 37242 6361
rect 37186 6287 37242 6296
rect 38384 6316 38436 6322
rect 34796 6248 34848 6254
rect 34796 6190 34848 6196
rect 34808 480 34836 6190
rect 35990 3496 36046 3505
rect 35990 3431 36046 3440
rect 36004 480 36032 3431
rect 37200 480 37228 6287
rect 38384 6258 38436 6264
rect 38396 480 38424 6258
rect 39592 480 39620 20334
rect 40696 480 40724 20470
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 41892 480 41920 3470
rect 43088 480 43116 22578
rect 43272 20602 43300 22100
rect 43260 20596 43312 20602
rect 43260 20538 43312 20544
rect 45468 20120 45520 20126
rect 45468 20062 45520 20068
rect 44272 5432 44324 5438
rect 44272 5374 44324 5380
rect 44284 480 44312 5374
rect 45480 480 45508 20062
rect 46676 480 46704 22578
rect 52552 22024 52604 22030
rect 52552 21966 52604 21972
rect 47860 21412 47912 21418
rect 47860 21354 47912 21360
rect 47872 480 47900 21354
rect 48964 5024 49016 5030
rect 48964 4966 49016 4972
rect 48976 480 49004 4966
rect 51356 3596 51408 3602
rect 51356 3538 51408 3544
rect 50160 3392 50212 3398
rect 50160 3334 50212 3340
rect 50172 480 50200 3334
rect 51368 480 51396 3538
rect 52564 480 52592 21966
rect 58440 21956 58492 21962
rect 58440 21898 58492 21904
rect 56048 6384 56100 6390
rect 56048 6326 56100 6332
rect 54942 4856 54998 4865
rect 54942 4791 54998 4800
rect 53748 3664 53800 3670
rect 53748 3606 53800 3612
rect 53760 480 53788 3606
rect 54956 480 54984 4791
rect 56060 480 56088 6326
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 57256 480 57284 3538
rect 58452 480 58480 21898
rect 59636 21888 59688 21894
rect 59636 21830 59688 21836
rect 59648 480 59676 21830
rect 65168 20262 65196 22100
rect 85592 22086 86434 22114
rect 65524 21820 65576 21826
rect 65524 21762 65576 21768
rect 65156 20256 65208 20262
rect 65156 20198 65208 20204
rect 64328 19984 64380 19990
rect 64328 19926 64380 19932
rect 63224 6452 63276 6458
rect 63224 6394 63276 6400
rect 62028 4140 62080 4146
rect 62028 4082 62080 4088
rect 60832 3664 60884 3670
rect 60832 3606 60884 3612
rect 60844 480 60872 3606
rect 62040 480 62068 4082
rect 63236 480 63264 6394
rect 64340 480 64368 19926
rect 65536 480 65564 21762
rect 73804 21752 73856 21758
rect 73804 21694 73856 21700
rect 70308 19780 70360 19786
rect 70308 19722 70360 19728
rect 66720 6520 66772 6526
rect 66720 6462 66772 6468
rect 66732 480 66760 6462
rect 69112 4956 69164 4962
rect 69112 4898 69164 4904
rect 67914 3632 67970 3641
rect 67914 3567 67970 3576
rect 67928 480 67956 3567
rect 69124 480 69152 4898
rect 70320 480 70348 19722
rect 72608 4956 72660 4962
rect 72608 4898 72660 4904
rect 71504 4072 71556 4078
rect 71504 4014 71556 4020
rect 71516 480 71544 4014
rect 72620 480 72648 4898
rect 73816 480 73844 21694
rect 84476 21684 84528 21690
rect 84476 21626 84528 21632
rect 82176 20596 82228 20602
rect 82176 20538 82228 20544
rect 78588 20460 78640 20466
rect 78588 20402 78640 20408
rect 76196 6860 76248 6866
rect 76196 6802 76248 6808
rect 75000 4004 75052 4010
rect 75000 3946 75052 3952
rect 75012 480 75040 3946
rect 76208 480 76236 6802
rect 77392 6520 77444 6526
rect 77392 6462 77444 6468
rect 77404 480 77432 6462
rect 78600 480 78628 20402
rect 80888 5024 80940 5030
rect 79690 4992 79746 5001
rect 80888 4966 80940 4972
rect 79690 4927 79746 4936
rect 79704 480 79732 4927
rect 80900 480 80928 4966
rect 82188 3874 82216 20538
rect 83280 5228 83332 5234
rect 83280 5170 83332 5176
rect 82084 3868 82136 3874
rect 82084 3810 82136 3816
rect 82176 3868 82228 3874
rect 82176 3810 82228 3816
rect 82096 480 82124 3810
rect 83292 480 83320 5170
rect 84488 480 84516 21626
rect 85592 3942 85620 22086
rect 86868 21616 86920 21622
rect 86868 21558 86920 21564
rect 85580 3936 85632 3942
rect 85580 3878 85632 3884
rect 85672 3800 85724 3806
rect 85672 3742 85724 3748
rect 85684 480 85712 3742
rect 86880 480 86908 21558
rect 89168 21548 89220 21554
rect 89168 21490 89220 21496
rect 87972 6588 88024 6594
rect 87972 6530 88024 6536
rect 87984 480 88012 6530
rect 89180 480 89208 21490
rect 90364 21480 90416 21486
rect 90364 21422 90416 21428
rect 90376 480 90404 21422
rect 98644 20256 98696 20262
rect 98644 20198 98696 20204
rect 93952 6792 94004 6798
rect 93952 6734 94004 6740
rect 92756 5092 92808 5098
rect 92756 5034 92808 5040
rect 91558 3768 91614 3777
rect 91558 3703 91614 3712
rect 91572 480 91600 3703
rect 92768 480 92796 5034
rect 93964 480 93992 6734
rect 97448 5228 97500 5234
rect 97448 5170 97500 5176
rect 96252 3732 96304 3738
rect 96252 3674 96304 3680
rect 95146 3224 95202 3233
rect 95146 3159 95202 3168
rect 95160 480 95188 3159
rect 96264 480 96292 3674
rect 97460 480 97488 5170
rect 98656 480 98684 20198
rect 102232 19916 102284 19922
rect 102232 19858 102284 19864
rect 101034 4992 101090 5001
rect 101034 4927 101090 4936
rect 99840 3800 99892 3806
rect 99840 3742 99892 3748
rect 99852 480 99880 3742
rect 101048 480 101076 4927
rect 102244 480 102272 19858
rect 108316 19378 108344 22100
rect 110510 21312 110566 21321
rect 110510 21247 110566 21256
rect 107016 19372 107068 19378
rect 107016 19314 107068 19320
rect 108304 19372 108356 19378
rect 108304 19314 108356 19320
rect 104532 5092 104584 5098
rect 104532 5034 104584 5040
rect 103336 3868 103388 3874
rect 103336 3810 103388 3816
rect 103348 480 103376 3810
rect 104544 480 104572 5034
rect 105728 3868 105780 3874
rect 105728 3810 105780 3816
rect 105740 480 105768 3810
rect 107028 3806 107056 19314
rect 108120 5296 108172 5302
rect 108120 5238 108172 5244
rect 107016 3800 107068 3806
rect 107016 3742 107068 3748
rect 106924 3732 106976 3738
rect 106924 3674 106976 3680
rect 106936 480 106964 3674
rect 108132 480 108160 5238
rect 109314 4040 109370 4049
rect 109314 3975 109370 3984
rect 109328 480 109356 3975
rect 110524 480 110552 21247
rect 114008 20596 114060 20602
rect 114008 20538 114060 20544
rect 112812 5364 112864 5370
rect 112812 5306 112864 5312
rect 111616 5296 111668 5302
rect 111616 5238 111668 5244
rect 111628 480 111656 5238
rect 112824 480 112852 5306
rect 114020 480 114048 20538
rect 129568 19854 129596 22100
rect 150452 22086 151478 22114
rect 129556 19848 129608 19854
rect 129556 19790 129608 19796
rect 150452 6866 150480 22086
rect 172716 19786 172744 22100
rect 172704 19780 172756 19786
rect 172704 19722 172756 19728
rect 150440 6860 150492 6866
rect 150440 6802 150492 6808
rect 194612 6798 194640 22100
rect 215864 20670 215892 22100
rect 215852 20664 215904 20670
rect 215852 20606 215904 20612
rect 237760 20534 237788 22100
rect 237748 20528 237800 20534
rect 237748 20470 237800 20476
rect 259012 19922 259040 22100
rect 280172 22086 280922 22114
rect 259000 19916 259052 19922
rect 259000 19858 259052 19864
rect 194600 6792 194652 6798
rect 194600 6734 194652 6740
rect 115204 6724 115256 6730
rect 115204 6666 115256 6672
rect 115216 480 115244 6666
rect 116400 6656 116452 6662
rect 116400 6598 116452 6604
rect 116412 480 116440 6598
rect 280172 5302 280200 22086
rect 302160 20602 302188 22100
rect 302148 20596 302200 20602
rect 302148 20538 302200 20544
rect 324056 20466 324084 22100
rect 324044 20460 324096 20466
rect 324044 20402 324096 20408
rect 345308 20398 345336 22100
rect 367112 22086 367218 22114
rect 345296 20392 345348 20398
rect 345296 20334 345348 20340
rect 367112 6730 367140 22086
rect 388456 20330 388484 22100
rect 388444 20324 388496 20330
rect 388444 20266 388496 20272
rect 410352 20194 410380 22100
rect 410340 20188 410392 20194
rect 410340 20130 410392 20136
rect 431604 20058 431632 22100
rect 453500 20126 453528 22100
rect 474752 20262 474780 22100
rect 495452 22086 496662 22114
rect 474740 20256 474792 20262
rect 474740 20198 474792 20204
rect 453488 20120 453540 20126
rect 453488 20062 453540 20068
rect 431592 20052 431644 20058
rect 431592 19994 431644 20000
rect 367100 6724 367152 6730
rect 367100 6666 367152 6672
rect 280160 5296 280212 5302
rect 122286 5264 122342 5273
rect 118620 5222 118832 5250
rect 118620 5166 118648 5222
rect 118608 5160 118660 5166
rect 118608 5102 118660 5108
rect 118700 5160 118752 5166
rect 118700 5102 118752 5108
rect 118712 3874 118740 5102
rect 118700 3868 118752 3874
rect 118700 3810 118752 3816
rect 117596 3800 117648 3806
rect 117596 3742 117648 3748
rect 117608 480 117636 3742
rect 118804 480 118832 5222
rect 280160 5238 280212 5244
rect 122286 5199 122342 5208
rect 119896 3936 119948 3942
rect 119896 3878 119948 3884
rect 121090 3904 121146 3913
rect 119908 480 119936 3878
rect 121090 3839 121146 3848
rect 121104 480 121132 3839
rect 122300 480 122328 5199
rect 123482 5128 123538 5137
rect 123482 5063 123538 5072
rect 123496 480 123524 5063
rect 495452 3942 495480 22086
rect 517900 19990 517928 22100
rect 539612 22086 539810 22114
rect 560312 22086 561062 22114
rect 517888 19984 517940 19990
rect 517888 19926 517940 19932
rect 539612 5234 539640 22086
rect 560312 6186 560340 22086
rect 561876 6458 561904 567559
rect 563072 499497 563100 679895
rect 563058 499488 563114 499497
rect 563058 499423 563114 499432
rect 563058 477048 563114 477057
rect 563058 476983 563114 476992
rect 561954 407824 562010 407833
rect 561954 407759 562010 407768
rect 561864 6452 561916 6458
rect 561864 6394 561916 6400
rect 560300 6180 560352 6186
rect 560300 6122 560352 6128
rect 539600 5228 539652 5234
rect 539600 5170 539652 5176
rect 561968 5030 561996 407759
rect 562046 385384 562102 385393
rect 562046 385319 562102 385328
rect 562060 6322 562088 385319
rect 562138 340368 562194 340377
rect 562138 340303 562194 340312
rect 562152 6390 562180 340303
rect 562230 294808 562286 294817
rect 562230 294743 562286 294752
rect 562140 6384 562192 6390
rect 562140 6326 562192 6332
rect 562048 6316 562100 6322
rect 562048 6258 562100 6264
rect 561956 5024 562008 5030
rect 561956 4966 562008 4972
rect 562244 4962 562272 294743
rect 562322 226128 562378 226137
rect 562322 226063 562378 226072
rect 562336 5098 562364 226063
rect 562414 135008 562470 135017
rect 562414 134943 562470 134952
rect 562428 6594 562456 134943
rect 562506 67008 562562 67017
rect 562506 66943 562562 66952
rect 562520 6662 562548 66943
rect 562598 43888 562654 43897
rect 562598 43823 562654 43832
rect 562508 6656 562560 6662
rect 562508 6598 562560 6604
rect 562416 6588 562468 6594
rect 562416 6530 562468 6536
rect 562612 6254 562640 43823
rect 562600 6248 562652 6254
rect 562600 6190 562652 6196
rect 562324 5092 562376 5098
rect 562324 5034 562376 5040
rect 562232 4956 562284 4962
rect 562232 4898 562284 4904
rect 495440 3936 495492 3942
rect 495440 3878 495492 3884
rect 124680 3868 124732 3874
rect 124680 3810 124732 3816
rect 124692 480 124720 3810
rect 563072 3670 563100 476983
rect 563150 431488 563206 431497
rect 563150 431423 563206 431432
rect 563164 3874 563192 431423
rect 563242 362808 563298 362817
rect 563242 362743 563298 362752
rect 563152 3868 563204 3874
rect 563152 3810 563204 3816
rect 563060 3664 563112 3670
rect 563060 3606 563112 3612
rect 563256 3369 563284 362743
rect 563334 317248 563390 317257
rect 563334 317183 563390 317192
rect 563348 3602 563376 317183
rect 563426 271688 563482 271697
rect 563426 271623 563482 271632
rect 563336 3596 563388 3602
rect 563336 3538 563388 3544
rect 563440 3534 563468 271623
rect 563518 249248 563574 249257
rect 563518 249183 563574 249192
rect 563532 5166 563560 249183
rect 563610 203688 563666 203697
rect 563610 203623 563666 203632
rect 563520 5160 563572 5166
rect 563520 5102 563572 5108
rect 563624 4826 563652 203623
rect 563702 180568 563758 180577
rect 563702 180503 563758 180512
rect 563716 4894 563744 180503
rect 563794 158128 563850 158137
rect 563794 158063 563850 158072
rect 563704 4888 563756 4894
rect 563704 4830 563756 4836
rect 563612 4820 563664 4826
rect 563612 4762 563664 4768
rect 563428 3528 563480 3534
rect 563428 3470 563480 3476
rect 563808 3466 563836 158063
rect 563886 112568 563942 112577
rect 563886 112503 563942 112512
rect 563900 6526 563928 112503
rect 563888 6520 563940 6526
rect 563888 6462 563940 6468
rect 564452 3806 564480 683198
rect 564532 683188 564584 683194
rect 564532 683130 564584 683136
rect 564440 3800 564492 3806
rect 564440 3742 564492 3748
rect 564544 3738 564572 683130
rect 564622 89448 564678 89457
rect 564622 89383 564678 89392
rect 564636 21418 564664 89383
rect 564624 21412 564676 21418
rect 564624 21354 564676 21360
rect 564532 3732 564584 3738
rect 564532 3674 564584 3680
rect 563796 3460 563848 3466
rect 563796 3402 563848 3408
rect 563242 3360 563298 3369
rect 563242 3295 563298 3304
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 4066 6160 4122 6216
rect 6458 3304 6514 3360
rect 17314 683440 17370 683496
rect 17682 683304 17738 683360
rect 18694 683576 18750 683632
rect 18602 363432 18658 363488
rect 19338 659912 19394 659968
rect 20166 614352 20222 614408
rect 19338 545672 19394 545728
rect 19338 500112 19394 500168
rect 21730 636792 21786 636848
rect 21638 591232 21694 591288
rect 20626 477672 20682 477728
rect 19706 454552 19762 454608
rect 20534 454552 20590 454608
rect 20534 408992 20590 409048
rect 20442 340992 20498 341048
rect 20350 317872 20406 317928
rect 20258 295432 20314 295488
rect 19338 272312 19394 272368
rect 20166 249872 20222 249928
rect 20074 204312 20130 204368
rect 19982 181192 20038 181248
rect 19522 135632 19578 135688
rect 19890 113192 19946 113248
rect 19798 67632 19854 67688
rect 19246 3168 19302 3224
rect 21546 386552 21602 386608
rect 21454 226752 21510 226808
rect 21362 158752 21418 158808
rect 21270 90072 21326 90128
rect 21178 44512 21234 44568
rect 345938 683848 345994 683904
rect 281538 683712 281594 683768
rect 324778 683168 324834 683224
rect 410982 683576 411038 683632
rect 432234 683440 432290 683496
rect 475382 683304 475438 683360
rect 21822 23432 21878 23488
rect 21730 3848 21786 3904
rect 367834 681264 367890 681320
rect 563058 679904 563114 679960
rect 561862 567568 561918 567624
rect 26514 22616 26570 22672
rect 33598 22616 33654 22672
rect 37186 6296 37242 6352
rect 35990 3440 36046 3496
rect 54942 4800 54998 4856
rect 67914 3576 67970 3632
rect 79690 4936 79746 4992
rect 91558 3712 91614 3768
rect 95146 3168 95202 3224
rect 101034 4936 101090 4992
rect 110510 21256 110566 21312
rect 109314 3984 109370 4040
rect 122286 5208 122342 5264
rect 121090 3848 121146 3904
rect 123482 5072 123538 5128
rect 563058 499432 563114 499488
rect 563058 476992 563114 477048
rect 561954 407768 562010 407824
rect 562046 385328 562102 385384
rect 562138 340312 562194 340368
rect 562230 294752 562286 294808
rect 562322 226072 562378 226128
rect 562414 134952 562470 135008
rect 562506 66952 562562 67008
rect 562598 43832 562654 43888
rect 563150 431432 563206 431488
rect 563242 362752 563298 362808
rect 563334 317192 563390 317248
rect 563426 271632 563482 271688
rect 563518 249192 563574 249248
rect 563610 203632 563666 203688
rect 563702 180512 563758 180568
rect 563794 158072 563850 158128
rect 563886 112512 563942 112568
rect 564622 89392 564678 89448
rect 563242 3304 563298 3360
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 21766 683844 21772 683908
rect 21836 683906 21842 683908
rect 345933 683906 345999 683909
rect 21836 683904 345999 683906
rect 21836 683848 345938 683904
rect 345994 683848 345999 683904
rect 21836 683846 345999 683848
rect 21836 683844 21842 683846
rect 345933 683843 345999 683846
rect 21950 683708 21956 683772
rect 22020 683770 22026 683772
rect 281533 683770 281599 683773
rect 22020 683768 281599 683770
rect 22020 683712 281538 683768
rect 281594 683712 281599 683768
rect 583520 683756 584960 683996
rect 22020 683710 281599 683712
rect 22020 683708 22026 683710
rect 281533 683707 281599 683710
rect 18689 683634 18755 683637
rect 410977 683634 411043 683637
rect 18689 683632 411043 683634
rect 18689 683576 18694 683632
rect 18750 683576 410982 683632
rect 411038 683576 411043 683632
rect 18689 683574 411043 683576
rect 18689 683571 18755 683574
rect 410977 683571 411043 683574
rect 17309 683498 17375 683501
rect 432229 683498 432295 683501
rect 17309 683496 432295 683498
rect 17309 683440 17314 683496
rect 17370 683440 432234 683496
rect 432290 683440 432295 683496
rect 17309 683438 432295 683440
rect 17309 683435 17375 683438
rect 432229 683435 432295 683438
rect 17677 683362 17743 683365
rect 475377 683362 475443 683365
rect 17677 683360 475443 683362
rect 17677 683304 17682 683360
rect 17738 683304 475382 683360
rect 475438 683304 475443 683360
rect 17677 683302 475443 683304
rect 17677 683299 17743 683302
rect 475377 683299 475443 683302
rect 324773 683226 324839 683229
rect 342110 683226 342116 683228
rect 324773 683224 342116 683226
rect 324773 683168 324778 683224
rect 324834 683168 342116 683224
rect 324773 683166 342116 683168
rect 324773 683163 324839 683166
rect 342110 683164 342116 683166
rect 342180 683164 342186 683228
rect 367829 681322 367895 681325
rect 354630 681320 367895 681322
rect 354630 681264 367834 681320
rect 367890 681264 367895 681320
rect 354630 681262 367895 681264
rect 21582 680444 21588 680508
rect 21652 680506 21658 680508
rect 354630 680506 354690 681262
rect 367829 681259 367895 681262
rect 21652 680446 354690 680506
rect 21652 680444 21658 680446
rect 342110 679900 342116 679964
rect 342180 679962 342186 679964
rect 563053 679962 563119 679965
rect 342180 679960 563119 679962
rect 342180 679904 563058 679960
rect 563114 679904 563119 679960
rect 342180 679902 563119 679904
rect 342180 679900 342186 679902
rect 563053 679899 563119 679902
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect 19333 659970 19399 659973
rect 19333 659968 22172 659970
rect 19333 659912 19338 659968
rect 19394 659912 22172 659968
rect 19333 659910 22172 659912
rect 19333 659907 19399 659910
rect 561622 659228 561628 659292
rect 561692 659228 561698 659292
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect 21725 636850 21791 636853
rect 21725 636848 22172 636850
rect 21725 636792 21730 636848
rect 21786 636792 22172 636848
rect 21725 636790 22172 636792
rect 21725 636787 21791 636790
rect 561806 636108 561812 636172
rect 561876 636108 561882 636172
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect 20161 614410 20227 614413
rect 20161 614408 22172 614410
rect 20161 614352 20166 614408
rect 20222 614352 22172 614408
rect 20161 614350 22172 614352
rect 20161 614347 20227 614350
rect 563094 613730 563100 613732
rect 561844 613670 563100 613730
rect 563094 613668 563100 613670
rect 563164 613668 563170 613732
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 21633 591290 21699 591293
rect 21633 591288 22172 591290
rect 21633 591232 21638 591288
rect 21694 591232 22172 591288
rect 21633 591230 22172 591232
rect 21633 591227 21699 591230
rect 583520 590868 584960 591108
rect 561814 590066 561874 590580
rect 561990 590066 561996 590068
rect 561814 590006 561996 590066
rect 561990 590004 561996 590006
rect 562060 590004 562066 590068
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect 20110 568788 20116 568852
rect 20180 568850 20186 568852
rect 20180 568790 22172 568850
rect 20180 568788 20186 568790
rect 561814 567629 561874 568140
rect 561814 567624 561923 567629
rect 561814 567568 561862 567624
rect 561918 567568 561923 567624
rect 561814 567566 561923 567568
rect 561857 567563 561923 567566
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect 19333 545730 19399 545733
rect 19333 545728 22172 545730
rect 19333 545672 19338 545728
rect 19394 545672 22172 545728
rect 19333 545670 22172 545672
rect 19333 545667 19399 545670
rect 562174 545050 562180 545052
rect 561844 544990 562180 545050
rect 562174 544988 562180 544990
rect 562244 544988 562250 545052
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect 19926 523228 19932 523292
rect 19996 523290 20002 523292
rect 19996 523230 22172 523290
rect 19996 523228 20002 523230
rect 563278 522610 563284 522612
rect 561844 522550 563284 522610
rect 563278 522548 563284 522550
rect 563348 522548 563354 522612
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 19333 500170 19399 500173
rect 19333 500168 22172 500170
rect 19333 500112 19338 500168
rect 19394 500112 22172 500168
rect 19333 500110 22172 500112
rect 19333 500107 19399 500110
rect 563053 499490 563119 499493
rect 561844 499488 563119 499490
rect 561844 499432 563058 499488
rect 563114 499432 563119 499488
rect 561844 499430 563119 499432
rect 563053 499427 563119 499430
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect 20621 477730 20687 477733
rect 20621 477728 22172 477730
rect 20621 477672 20626 477728
rect 20682 477672 22172 477728
rect 20621 477670 22172 477672
rect 20621 477667 20687 477670
rect 563053 477050 563119 477053
rect 561844 477048 563119 477050
rect 561844 476992 563058 477048
rect 563114 476992 563119 477048
rect 561844 476990 563119 476992
rect 563053 476987 563119 476990
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect 19701 454610 19767 454613
rect 20529 454610 20595 454613
rect 19701 454608 22172 454610
rect 19701 454552 19706 454608
rect 19762 454552 20534 454608
rect 20590 454552 22172 454608
rect 19701 454550 22172 454552
rect 19701 454547 19767 454550
rect 20529 454547 20595 454550
rect 563462 453930 563468 453932
rect 561844 453870 563468 453930
rect 563462 453868 563468 453870
rect 563532 453868 563538 453932
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 19742 432108 19748 432172
rect 19812 432170 19818 432172
rect 19812 432110 22172 432170
rect 19812 432108 19818 432110
rect 563145 431490 563211 431493
rect 561844 431488 563211 431490
rect 561844 431432 563150 431488
rect 563206 431432 563211 431488
rect 583520 431476 584960 431716
rect 561844 431430 563211 431432
rect 563145 431427 563211 431430
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 20529 409050 20595 409053
rect 20529 409048 22172 409050
rect 20529 408992 20534 409048
rect 20590 408992 22172 409048
rect 20529 408990 22172 408992
rect 20529 408987 20595 408990
rect 561814 407826 561874 408340
rect 561949 407826 562015 407829
rect 561814 407824 562015 407826
rect 561814 407768 561954 407824
rect 562010 407768 562015 407824
rect 561814 407766 562015 407768
rect 561949 407763 562015 407766
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect 21541 386610 21607 386613
rect 21541 386608 22172 386610
rect 21541 386552 21546 386608
rect 21602 386552 22172 386608
rect 21541 386550 22172 386552
rect 21541 386547 21607 386550
rect 561814 385386 561874 385900
rect 562041 385386 562107 385389
rect 561814 385384 562107 385386
rect 561814 385328 562046 385384
rect 562102 385328 562107 385384
rect 561814 385326 562107 385328
rect 562041 385323 562107 385326
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect 18597 363490 18663 363493
rect 18597 363488 22172 363490
rect 18597 363432 18602 363488
rect 18658 363432 22172 363488
rect 18597 363430 22172 363432
rect 18597 363427 18663 363430
rect 563237 362810 563303 362813
rect 561844 362808 563303 362810
rect 561844 362752 563242 362808
rect 563298 362752 563303 362808
rect 561844 362750 563303 362752
rect 563237 362747 563303 362750
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 20437 341050 20503 341053
rect 20437 341048 22172 341050
rect 20437 340992 20442 341048
rect 20498 340992 22172 341048
rect 20437 340990 22172 340992
rect 20437 340987 20503 340990
rect 562133 340370 562199 340373
rect 561844 340368 562199 340370
rect 561844 340312 562138 340368
rect 562194 340312 562199 340368
rect 561844 340310 562199 340312
rect 562133 340307 562199 340310
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 20345 317930 20411 317933
rect 20345 317928 22172 317930
rect 20345 317872 20350 317928
rect 20406 317872 22172 317928
rect 20345 317870 22172 317872
rect 20345 317867 20411 317870
rect 563329 317250 563395 317253
rect 561844 317248 563395 317250
rect 561844 317192 563334 317248
rect 563390 317192 563395 317248
rect 561844 317190 563395 317192
rect 563329 317187 563395 317190
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect 20253 295490 20319 295493
rect 20253 295488 22172 295490
rect 20253 295432 20258 295488
rect 20314 295432 22172 295488
rect 20253 295430 22172 295432
rect 20253 295427 20319 295430
rect 562225 294810 562291 294813
rect 561844 294808 562291 294810
rect 561844 294752 562230 294808
rect 562286 294752 562291 294808
rect 561844 294750 562291 294752
rect 562225 294747 562291 294750
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 19333 272370 19399 272373
rect 19333 272368 22172 272370
rect 19333 272312 19338 272368
rect 19394 272312 22172 272368
rect 19333 272310 22172 272312
rect 19333 272307 19399 272310
rect 583520 272084 584960 272324
rect 563421 271690 563487 271693
rect 561844 271688 563487 271690
rect 561844 271632 563426 271688
rect 563482 271632 563487 271688
rect 561844 271630 563487 271632
rect 563421 271627 563487 271630
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 20161 249930 20227 249933
rect 20161 249928 22172 249930
rect 20161 249872 20166 249928
rect 20222 249872 22172 249928
rect 20161 249870 22172 249872
rect 20161 249867 20227 249870
rect 563513 249250 563579 249253
rect 561844 249248 563579 249250
rect 561844 249192 563518 249248
rect 563574 249192 563579 249248
rect 561844 249190 563579 249192
rect 563513 249187 563579 249190
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 21449 226810 21515 226813
rect 21449 226808 22172 226810
rect 21449 226752 21454 226808
rect 21510 226752 22172 226808
rect 21449 226750 22172 226752
rect 21449 226747 21515 226750
rect 562317 226130 562383 226133
rect 561844 226128 562383 226130
rect 561844 226072 562322 226128
rect 562378 226072 562383 226128
rect 561844 226070 562383 226072
rect 562317 226067 562383 226070
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect 20069 204370 20135 204373
rect 20069 204368 22172 204370
rect 20069 204312 20074 204368
rect 20130 204312 22172 204368
rect 20069 204310 22172 204312
rect 20069 204307 20135 204310
rect 563605 203690 563671 203693
rect 561844 203688 563671 203690
rect 561844 203632 563610 203688
rect 563666 203632 563671 203688
rect 561844 203630 563671 203632
rect 563605 203627 563671 203630
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 19977 181250 20043 181253
rect 19977 181248 22172 181250
rect 19977 181192 19982 181248
rect 20038 181192 22172 181248
rect 19977 181190 22172 181192
rect 19977 181187 20043 181190
rect 563697 180570 563763 180573
rect 561844 180568 563763 180570
rect 561844 180512 563702 180568
rect 563758 180512 563763 180568
rect 561844 180510 563763 180512
rect 563697 180507 563763 180510
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 21357 158810 21423 158813
rect 21357 158808 22172 158810
rect 21357 158752 21362 158808
rect 21418 158752 22172 158808
rect 21357 158750 22172 158752
rect 21357 158747 21423 158750
rect 563789 158130 563855 158133
rect 561844 158128 563855 158130
rect 561844 158072 563794 158128
rect 563850 158072 563855 158128
rect 561844 158070 563855 158072
rect 563789 158067 563855 158070
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 19517 135690 19583 135693
rect 19517 135688 22172 135690
rect 19517 135632 19522 135688
rect 19578 135632 22172 135688
rect 19517 135630 22172 135632
rect 19517 135627 19583 135630
rect 562409 135010 562475 135013
rect 561844 135008 562475 135010
rect 561844 134952 562414 135008
rect 562470 134952 562475 135008
rect 561844 134950 562475 134952
rect 562409 134947 562475 134950
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 19885 113250 19951 113253
rect 19885 113248 22172 113250
rect 19885 113192 19890 113248
rect 19946 113192 22172 113248
rect 19885 113190 22172 113192
rect 19885 113187 19951 113190
rect 583520 112692 584960 112932
rect 563881 112570 563947 112573
rect 561844 112568 563947 112570
rect 561844 112512 563886 112568
rect 563942 112512 563947 112568
rect 561844 112510 563947 112512
rect 563881 112507 563947 112510
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 21265 90130 21331 90133
rect 21265 90128 22172 90130
rect 21265 90072 21270 90128
rect 21326 90072 22172 90128
rect 21265 90070 22172 90072
rect 21265 90067 21331 90070
rect 564617 89450 564683 89453
rect 561844 89448 564683 89450
rect 561844 89392 564622 89448
rect 564678 89392 564683 89448
rect 561844 89390 564683 89392
rect 564617 89387 564683 89390
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 19793 67690 19859 67693
rect 19793 67688 22172 67690
rect 19793 67632 19798 67688
rect 19854 67632 22172 67688
rect 19793 67630 22172 67632
rect 19793 67627 19859 67630
rect 562501 67010 562567 67013
rect 561844 67008 562567 67010
rect 561844 66952 562506 67008
rect 562562 66952 562567 67008
rect 561844 66950 562567 66952
rect 562501 66947 562567 66950
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 21173 44570 21239 44573
rect 21173 44568 22172 44570
rect 21173 44512 21178 44568
rect 21234 44512 22172 44568
rect 21173 44510 22172 44512
rect 21173 44507 21239 44510
rect 562593 43890 562659 43893
rect 561844 43888 562659 43890
rect 561844 43832 562598 43888
rect 562654 43832 562659 43888
rect 561844 43830 562659 43832
rect 562593 43827 562659 43830
rect 21582 42876 21588 42940
rect 21652 42938 21658 42940
rect 22502 42938 22508 42940
rect 21652 42878 22508 42938
rect 21652 42876 21658 42878
rect 22502 42876 22508 42878
rect 22572 42876 22578 42940
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 21817 23490 21883 23493
rect 23790 23490 23796 23492
rect 21817 23488 23796 23490
rect 21817 23432 21822 23488
rect 21878 23432 23796 23488
rect 21817 23430 23796 23432
rect 21817 23427 21883 23430
rect 23790 23428 23796 23430
rect 23860 23428 23866 23492
rect 21766 22748 21772 22812
rect 21836 22810 21842 22812
rect 21836 22750 29930 22810
rect 21836 22748 21842 22750
rect 21950 22612 21956 22676
rect 22020 22674 22026 22676
rect 26509 22674 26575 22677
rect 22020 22672 26575 22674
rect 22020 22616 26514 22672
rect 26570 22616 26575 22672
rect 22020 22614 26575 22616
rect 29870 22674 29930 22750
rect 33593 22674 33659 22677
rect 29870 22672 33659 22674
rect 29870 22616 33598 22672
rect 33654 22616 33659 22672
rect 29870 22614 33659 22616
rect 22020 22612 22026 22614
rect 26509 22611 26575 22614
rect 33593 22611 33659 22614
rect 22686 21252 22692 21316
rect 22756 21314 22762 21316
rect 110505 21314 110571 21317
rect 22756 21312 110571 21314
rect 22756 21256 110510 21312
rect 110566 21256 110571 21312
rect 22756 21254 110571 21256
rect 22756 21252 22762 21254
rect 110505 21251 110571 21254
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 37181 6354 37247 6357
rect 562174 6354 562180 6356
rect 37181 6352 562180 6354
rect 37181 6296 37186 6352
rect 37242 6296 562180 6352
rect 37181 6294 562180 6296
rect 37181 6291 37247 6294
rect 562174 6292 562180 6294
rect 562244 6292 562250 6356
rect 4061 6218 4127 6221
rect 563094 6218 563100 6220
rect 4061 6216 563100 6218
rect 4061 6160 4066 6216
rect 4122 6160 563100 6216
rect 4061 6158 563100 6160
rect 4061 6155 4127 6158
rect 563094 6156 563100 6158
rect 563164 6156 563170 6220
rect 19742 5204 19748 5268
rect 19812 5266 19818 5268
rect 122281 5266 122347 5269
rect 19812 5264 122347 5266
rect 19812 5208 122286 5264
rect 122342 5208 122347 5264
rect 19812 5206 122347 5208
rect 19812 5204 19818 5206
rect 122281 5203 122347 5206
rect 20110 5068 20116 5132
rect 20180 5130 20186 5132
rect 123477 5130 123543 5133
rect 20180 5128 123543 5130
rect 20180 5072 123482 5128
rect 123538 5072 123543 5128
rect 20180 5070 123543 5072
rect 20180 5068 20186 5070
rect 123477 5067 123543 5070
rect 19926 4932 19932 4996
rect 19996 4994 20002 4996
rect 79685 4994 79751 4997
rect 19996 4992 79751 4994
rect 19996 4936 79690 4992
rect 79746 4936 79751 4992
rect 19996 4934 79751 4936
rect 19996 4932 20002 4934
rect 79685 4931 79751 4934
rect 101029 4994 101095 4997
rect 561622 4994 561628 4996
rect 101029 4992 561628 4994
rect 101029 4936 101034 4992
rect 101090 4936 561628 4992
rect 101029 4934 561628 4936
rect 101029 4931 101095 4934
rect 561622 4932 561628 4934
rect 561692 4932 561698 4996
rect 54937 4858 55003 4861
rect 561990 4858 561996 4860
rect 54937 4856 561996 4858
rect 54937 4800 54942 4856
rect 54998 4800 561996 4856
rect 54937 4798 561996 4800
rect 54937 4795 55003 4798
rect 561990 4796 561996 4798
rect 562060 4796 562066 4860
rect 23790 3980 23796 4044
rect 23860 4042 23866 4044
rect 109309 4042 109375 4045
rect 23860 4040 109375 4042
rect 23860 3984 109314 4040
rect 109370 3984 109375 4040
rect 23860 3982 109375 3984
rect 23860 3980 23866 3982
rect 109309 3979 109375 3982
rect 21725 3906 21791 3909
rect 121085 3906 121151 3909
rect 21725 3904 121151 3906
rect 21725 3848 21730 3904
rect 21786 3848 121090 3904
rect 121146 3848 121151 3904
rect 21725 3846 121151 3848
rect 21725 3843 21791 3846
rect 121085 3843 121151 3846
rect 91553 3770 91619 3773
rect 561806 3770 561812 3772
rect 91553 3768 561812 3770
rect 91553 3712 91558 3768
rect 91614 3712 561812 3768
rect 91553 3710 561812 3712
rect 91553 3707 91619 3710
rect 561806 3708 561812 3710
rect 561876 3708 561882 3772
rect 67909 3634 67975 3637
rect 563278 3634 563284 3636
rect 67909 3632 563284 3634
rect 67909 3576 67914 3632
rect 67970 3576 563284 3632
rect 67909 3574 563284 3576
rect 67909 3571 67975 3574
rect 563278 3572 563284 3574
rect 563348 3572 563354 3636
rect 35985 3498 36051 3501
rect 563462 3498 563468 3500
rect 35985 3496 563468 3498
rect 35985 3440 35990 3496
rect 36046 3440 563468 3496
rect 35985 3438 563468 3440
rect 35985 3435 36051 3438
rect 563462 3436 563468 3438
rect 563532 3436 563538 3500
rect 6453 3362 6519 3365
rect 563237 3362 563303 3365
rect 6453 3360 563303 3362
rect 6453 3304 6458 3360
rect 6514 3304 563242 3360
rect 563298 3304 563303 3360
rect 6453 3302 563303 3304
rect 6453 3299 6519 3302
rect 563237 3299 563303 3302
rect 19241 3226 19307 3229
rect 95141 3226 95207 3229
rect 19241 3224 95207 3226
rect 19241 3168 19246 3224
rect 19302 3168 95146 3224
rect 95202 3168 95207 3224
rect 19241 3166 95207 3168
rect 19241 3163 19307 3166
rect 95141 3163 95207 3166
<< via3 >>
rect 21772 683844 21836 683908
rect 21956 683708 22020 683772
rect 342116 683164 342180 683228
rect 21588 680444 21652 680508
rect 342116 679900 342180 679964
rect 561628 659228 561692 659292
rect 561812 636108 561876 636172
rect 563100 613668 563164 613732
rect 561996 590004 562060 590068
rect 20116 568788 20180 568852
rect 562180 544988 562244 545052
rect 19932 523228 19996 523292
rect 563284 522548 563348 522612
rect 563468 453868 563532 453932
rect 19748 432108 19812 432172
rect 21588 42876 21652 42940
rect 22508 42876 22572 42940
rect 23796 23428 23860 23492
rect 21772 22748 21836 22812
rect 21956 22612 22020 22676
rect 22692 21252 22756 21316
rect 562180 6292 562244 6356
rect 563100 6156 563164 6220
rect 19748 5204 19812 5268
rect 20116 5068 20180 5132
rect 19932 4932 19996 4996
rect 561628 4932 561692 4996
rect 561996 4796 562060 4860
rect 23796 3980 23860 4044
rect 561812 3708 561876 3772
rect 563284 3572 563348 3636
rect 563468 3436 563532 3500
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 21771 683908 21837 683909
rect 21771 683844 21772 683908
rect 21836 683844 21837 683908
rect 21771 683843 21837 683844
rect 21587 680508 21653 680509
rect 21587 680444 21588 680508
rect 21652 680444 21653 680508
rect 21587 680443 21653 680444
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20115 568852 20181 568853
rect 20115 568788 20116 568852
rect 20180 568788 20181 568852
rect 20115 568787 20181 568788
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 19931 523292 19997 523293
rect 19931 523228 19932 523292
rect 19996 523228 19997 523292
rect 19931 523227 19997 523228
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 19747 432172 19813 432173
rect 19747 432108 19748 432172
rect 19812 432108 19813 432172
rect 19747 432107 19813 432108
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 19750 5269 19810 432107
rect 19747 5268 19813 5269
rect 19747 5204 19748 5268
rect 19812 5204 19813 5268
rect 19747 5203 19813 5204
rect 19934 4997 19994 523227
rect 20118 5133 20178 568787
rect 20394 562054 21014 597498
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 21590 42941 21650 680443
rect 21587 42940 21653 42941
rect 21587 42876 21588 42940
rect 21652 42876 21653 42940
rect 21587 42875 21653 42876
rect 21774 22813 21834 683843
rect 21955 683772 22021 683773
rect 21955 683708 21956 683772
rect 22020 683708 22021 683772
rect 21955 683707 22021 683708
rect 21771 22812 21837 22813
rect 21771 22748 21772 22812
rect 21836 22748 21837 22812
rect 21771 22747 21837 22748
rect 21958 22677 22018 683707
rect 24114 673774 24734 710042
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 681449 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 681804 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 681449 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 681449 49574 698058
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 681449 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 681449 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 681449 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 681449 85574 698058
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 681449 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 681449 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 681449 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 681449 121574 698058
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 681449 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 681449 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 681449 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 681449 157574 698058
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 681449 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 681449 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 681449 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 681449 193574 698058
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 681449 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 681449 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 681804 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 681449 229574 698058
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 681449 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 681449 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 681449 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 681449 265574 698058
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 681449 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 681449 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 681449 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 681449 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 681449 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 681449 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 681804 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 681449 337574 698058
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 342115 683228 342181 683229
rect 342115 683164 342116 683228
rect 342180 683164 342181 683228
rect 342115 683163 342181 683164
rect 342118 679965 342178 683163
rect 361794 681449 362414 686898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 681449 366134 690618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 681449 369854 694338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 681449 373574 698058
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 681449 398414 686898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 681449 402134 690618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 681449 405854 694338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 681449 409574 698058
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 681449 434414 686898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 681449 438134 690618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 681804 441854 694338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 681449 445574 698058
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 681449 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 681449 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 681449 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 681449 481574 698058
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 681449 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 681449 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 681449 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 681449 517574 698058
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 681449 542414 686898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 681449 546134 690618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 681449 549854 694338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 681449 553574 698058
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 342115 679964 342181 679965
rect 342115 679900 342116 679964
rect 342180 679900 342181 679964
rect 342115 679899 342181 679900
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 637774 24734 673218
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 41568 655174 41888 655206
rect 41568 654938 41610 655174
rect 41846 654938 41888 655174
rect 41568 654854 41888 654938
rect 41568 654618 41610 654854
rect 41846 654618 41888 654854
rect 41568 654586 41888 654618
rect 72288 655174 72608 655206
rect 72288 654938 72330 655174
rect 72566 654938 72608 655174
rect 72288 654854 72608 654938
rect 72288 654618 72330 654854
rect 72566 654618 72608 654854
rect 72288 654586 72608 654618
rect 103008 655174 103328 655206
rect 103008 654938 103050 655174
rect 103286 654938 103328 655174
rect 103008 654854 103328 654938
rect 103008 654618 103050 654854
rect 103286 654618 103328 654854
rect 103008 654586 103328 654618
rect 133728 655174 134048 655206
rect 133728 654938 133770 655174
rect 134006 654938 134048 655174
rect 133728 654854 134048 654938
rect 133728 654618 133770 654854
rect 134006 654618 134048 654854
rect 133728 654586 134048 654618
rect 164448 655174 164768 655206
rect 164448 654938 164490 655174
rect 164726 654938 164768 655174
rect 164448 654854 164768 654938
rect 164448 654618 164490 654854
rect 164726 654618 164768 654854
rect 164448 654586 164768 654618
rect 195168 655174 195488 655206
rect 195168 654938 195210 655174
rect 195446 654938 195488 655174
rect 195168 654854 195488 654938
rect 195168 654618 195210 654854
rect 195446 654618 195488 654854
rect 195168 654586 195488 654618
rect 225888 655174 226208 655206
rect 225888 654938 225930 655174
rect 226166 654938 226208 655174
rect 225888 654854 226208 654938
rect 225888 654618 225930 654854
rect 226166 654618 226208 654854
rect 225888 654586 226208 654618
rect 256608 655174 256928 655206
rect 256608 654938 256650 655174
rect 256886 654938 256928 655174
rect 256608 654854 256928 654938
rect 256608 654618 256650 654854
rect 256886 654618 256928 654854
rect 256608 654586 256928 654618
rect 287328 655174 287648 655206
rect 287328 654938 287370 655174
rect 287606 654938 287648 655174
rect 287328 654854 287648 654938
rect 287328 654618 287370 654854
rect 287606 654618 287648 654854
rect 287328 654586 287648 654618
rect 318048 655174 318368 655206
rect 318048 654938 318090 655174
rect 318326 654938 318368 655174
rect 318048 654854 318368 654938
rect 318048 654618 318090 654854
rect 318326 654618 318368 654854
rect 318048 654586 318368 654618
rect 348768 655174 349088 655206
rect 348768 654938 348810 655174
rect 349046 654938 349088 655174
rect 348768 654854 349088 654938
rect 348768 654618 348810 654854
rect 349046 654618 349088 654854
rect 348768 654586 349088 654618
rect 379488 655174 379808 655206
rect 379488 654938 379530 655174
rect 379766 654938 379808 655174
rect 379488 654854 379808 654938
rect 379488 654618 379530 654854
rect 379766 654618 379808 654854
rect 379488 654586 379808 654618
rect 410208 655174 410528 655206
rect 410208 654938 410250 655174
rect 410486 654938 410528 655174
rect 410208 654854 410528 654938
rect 410208 654618 410250 654854
rect 410486 654618 410528 654854
rect 410208 654586 410528 654618
rect 440928 655174 441248 655206
rect 440928 654938 440970 655174
rect 441206 654938 441248 655174
rect 440928 654854 441248 654938
rect 440928 654618 440970 654854
rect 441206 654618 441248 654854
rect 440928 654586 441248 654618
rect 471648 655174 471968 655206
rect 471648 654938 471690 655174
rect 471926 654938 471968 655174
rect 471648 654854 471968 654938
rect 471648 654618 471690 654854
rect 471926 654618 471968 654854
rect 471648 654586 471968 654618
rect 502368 655174 502688 655206
rect 502368 654938 502410 655174
rect 502646 654938 502688 655174
rect 502368 654854 502688 654938
rect 502368 654618 502410 654854
rect 502646 654618 502688 654854
rect 502368 654586 502688 654618
rect 533088 655174 533408 655206
rect 533088 654938 533130 655174
rect 533366 654938 533408 655174
rect 533088 654854 533408 654938
rect 533088 654618 533130 654854
rect 533366 654618 533408 654854
rect 533088 654586 533408 654618
rect 26208 651454 26528 651486
rect 26208 651218 26250 651454
rect 26486 651218 26528 651454
rect 26208 651134 26528 651218
rect 26208 650898 26250 651134
rect 26486 650898 26528 651134
rect 26208 650866 26528 650898
rect 56928 651454 57248 651486
rect 56928 651218 56970 651454
rect 57206 651218 57248 651454
rect 56928 651134 57248 651218
rect 56928 650898 56970 651134
rect 57206 650898 57248 651134
rect 56928 650866 57248 650898
rect 87648 651454 87968 651486
rect 87648 651218 87690 651454
rect 87926 651218 87968 651454
rect 87648 651134 87968 651218
rect 87648 650898 87690 651134
rect 87926 650898 87968 651134
rect 87648 650866 87968 650898
rect 118368 651454 118688 651486
rect 118368 651218 118410 651454
rect 118646 651218 118688 651454
rect 118368 651134 118688 651218
rect 118368 650898 118410 651134
rect 118646 650898 118688 651134
rect 118368 650866 118688 650898
rect 149088 651454 149408 651486
rect 149088 651218 149130 651454
rect 149366 651218 149408 651454
rect 149088 651134 149408 651218
rect 149088 650898 149130 651134
rect 149366 650898 149408 651134
rect 149088 650866 149408 650898
rect 179808 651454 180128 651486
rect 179808 651218 179850 651454
rect 180086 651218 180128 651454
rect 179808 651134 180128 651218
rect 179808 650898 179850 651134
rect 180086 650898 180128 651134
rect 179808 650866 180128 650898
rect 210528 651454 210848 651486
rect 210528 651218 210570 651454
rect 210806 651218 210848 651454
rect 210528 651134 210848 651218
rect 210528 650898 210570 651134
rect 210806 650898 210848 651134
rect 210528 650866 210848 650898
rect 241248 651454 241568 651486
rect 241248 651218 241290 651454
rect 241526 651218 241568 651454
rect 241248 651134 241568 651218
rect 241248 650898 241290 651134
rect 241526 650898 241568 651134
rect 241248 650866 241568 650898
rect 271968 651454 272288 651486
rect 271968 651218 272010 651454
rect 272246 651218 272288 651454
rect 271968 651134 272288 651218
rect 271968 650898 272010 651134
rect 272246 650898 272288 651134
rect 271968 650866 272288 650898
rect 302688 651454 303008 651486
rect 302688 651218 302730 651454
rect 302966 651218 303008 651454
rect 302688 651134 303008 651218
rect 302688 650898 302730 651134
rect 302966 650898 303008 651134
rect 302688 650866 303008 650898
rect 333408 651454 333728 651486
rect 333408 651218 333450 651454
rect 333686 651218 333728 651454
rect 333408 651134 333728 651218
rect 333408 650898 333450 651134
rect 333686 650898 333728 651134
rect 333408 650866 333728 650898
rect 364128 651454 364448 651486
rect 364128 651218 364170 651454
rect 364406 651218 364448 651454
rect 364128 651134 364448 651218
rect 364128 650898 364170 651134
rect 364406 650898 364448 651134
rect 364128 650866 364448 650898
rect 394848 651454 395168 651486
rect 394848 651218 394890 651454
rect 395126 651218 395168 651454
rect 394848 651134 395168 651218
rect 394848 650898 394890 651134
rect 395126 650898 395168 651134
rect 394848 650866 395168 650898
rect 425568 651454 425888 651486
rect 425568 651218 425610 651454
rect 425846 651218 425888 651454
rect 425568 651134 425888 651218
rect 425568 650898 425610 651134
rect 425846 650898 425888 651134
rect 425568 650866 425888 650898
rect 456288 651454 456608 651486
rect 456288 651218 456330 651454
rect 456566 651218 456608 651454
rect 456288 651134 456608 651218
rect 456288 650898 456330 651134
rect 456566 650898 456608 651134
rect 456288 650866 456608 650898
rect 487008 651454 487328 651486
rect 487008 651218 487050 651454
rect 487286 651218 487328 651454
rect 487008 651134 487328 651218
rect 487008 650898 487050 651134
rect 487286 650898 487328 651134
rect 487008 650866 487328 650898
rect 517728 651454 518048 651486
rect 517728 651218 517770 651454
rect 518006 651218 518048 651454
rect 517728 651134 518048 651218
rect 517728 650898 517770 651134
rect 518006 650898 518048 651134
rect 517728 650866 518048 650898
rect 548448 651454 548768 651486
rect 548448 651218 548490 651454
rect 548726 651218 548768 651454
rect 548448 651134 548768 651218
rect 548448 650898 548490 651134
rect 548726 650898 548768 651134
rect 548448 650866 548768 650898
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 601774 24734 637218
rect 560394 634054 561014 669498
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 561627 659292 561693 659293
rect 561627 659228 561628 659292
rect 561692 659228 561693 659292
rect 561627 659227 561693 659228
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 41568 619174 41888 619206
rect 41568 618938 41610 619174
rect 41846 618938 41888 619174
rect 41568 618854 41888 618938
rect 41568 618618 41610 618854
rect 41846 618618 41888 618854
rect 41568 618586 41888 618618
rect 72288 619174 72608 619206
rect 72288 618938 72330 619174
rect 72566 618938 72608 619174
rect 72288 618854 72608 618938
rect 72288 618618 72330 618854
rect 72566 618618 72608 618854
rect 72288 618586 72608 618618
rect 103008 619174 103328 619206
rect 103008 618938 103050 619174
rect 103286 618938 103328 619174
rect 103008 618854 103328 618938
rect 103008 618618 103050 618854
rect 103286 618618 103328 618854
rect 103008 618586 103328 618618
rect 133728 619174 134048 619206
rect 133728 618938 133770 619174
rect 134006 618938 134048 619174
rect 133728 618854 134048 618938
rect 133728 618618 133770 618854
rect 134006 618618 134048 618854
rect 133728 618586 134048 618618
rect 164448 619174 164768 619206
rect 164448 618938 164490 619174
rect 164726 618938 164768 619174
rect 164448 618854 164768 618938
rect 164448 618618 164490 618854
rect 164726 618618 164768 618854
rect 164448 618586 164768 618618
rect 195168 619174 195488 619206
rect 195168 618938 195210 619174
rect 195446 618938 195488 619174
rect 195168 618854 195488 618938
rect 195168 618618 195210 618854
rect 195446 618618 195488 618854
rect 195168 618586 195488 618618
rect 225888 619174 226208 619206
rect 225888 618938 225930 619174
rect 226166 618938 226208 619174
rect 225888 618854 226208 618938
rect 225888 618618 225930 618854
rect 226166 618618 226208 618854
rect 225888 618586 226208 618618
rect 256608 619174 256928 619206
rect 256608 618938 256650 619174
rect 256886 618938 256928 619174
rect 256608 618854 256928 618938
rect 256608 618618 256650 618854
rect 256886 618618 256928 618854
rect 256608 618586 256928 618618
rect 287328 619174 287648 619206
rect 287328 618938 287370 619174
rect 287606 618938 287648 619174
rect 287328 618854 287648 618938
rect 287328 618618 287370 618854
rect 287606 618618 287648 618854
rect 287328 618586 287648 618618
rect 318048 619174 318368 619206
rect 318048 618938 318090 619174
rect 318326 618938 318368 619174
rect 318048 618854 318368 618938
rect 318048 618618 318090 618854
rect 318326 618618 318368 618854
rect 318048 618586 318368 618618
rect 348768 619174 349088 619206
rect 348768 618938 348810 619174
rect 349046 618938 349088 619174
rect 348768 618854 349088 618938
rect 348768 618618 348810 618854
rect 349046 618618 349088 618854
rect 348768 618586 349088 618618
rect 379488 619174 379808 619206
rect 379488 618938 379530 619174
rect 379766 618938 379808 619174
rect 379488 618854 379808 618938
rect 379488 618618 379530 618854
rect 379766 618618 379808 618854
rect 379488 618586 379808 618618
rect 410208 619174 410528 619206
rect 410208 618938 410250 619174
rect 410486 618938 410528 619174
rect 410208 618854 410528 618938
rect 410208 618618 410250 618854
rect 410486 618618 410528 618854
rect 410208 618586 410528 618618
rect 440928 619174 441248 619206
rect 440928 618938 440970 619174
rect 441206 618938 441248 619174
rect 440928 618854 441248 618938
rect 440928 618618 440970 618854
rect 441206 618618 441248 618854
rect 440928 618586 441248 618618
rect 471648 619174 471968 619206
rect 471648 618938 471690 619174
rect 471926 618938 471968 619174
rect 471648 618854 471968 618938
rect 471648 618618 471690 618854
rect 471926 618618 471968 618854
rect 471648 618586 471968 618618
rect 502368 619174 502688 619206
rect 502368 618938 502410 619174
rect 502646 618938 502688 619174
rect 502368 618854 502688 618938
rect 502368 618618 502410 618854
rect 502646 618618 502688 618854
rect 502368 618586 502688 618618
rect 533088 619174 533408 619206
rect 533088 618938 533130 619174
rect 533366 618938 533408 619174
rect 533088 618854 533408 618938
rect 533088 618618 533130 618854
rect 533366 618618 533408 618854
rect 533088 618586 533408 618618
rect 26208 615454 26528 615486
rect 26208 615218 26250 615454
rect 26486 615218 26528 615454
rect 26208 615134 26528 615218
rect 26208 614898 26250 615134
rect 26486 614898 26528 615134
rect 26208 614866 26528 614898
rect 56928 615454 57248 615486
rect 56928 615218 56970 615454
rect 57206 615218 57248 615454
rect 56928 615134 57248 615218
rect 56928 614898 56970 615134
rect 57206 614898 57248 615134
rect 56928 614866 57248 614898
rect 87648 615454 87968 615486
rect 87648 615218 87690 615454
rect 87926 615218 87968 615454
rect 87648 615134 87968 615218
rect 87648 614898 87690 615134
rect 87926 614898 87968 615134
rect 87648 614866 87968 614898
rect 118368 615454 118688 615486
rect 118368 615218 118410 615454
rect 118646 615218 118688 615454
rect 118368 615134 118688 615218
rect 118368 614898 118410 615134
rect 118646 614898 118688 615134
rect 118368 614866 118688 614898
rect 149088 615454 149408 615486
rect 149088 615218 149130 615454
rect 149366 615218 149408 615454
rect 149088 615134 149408 615218
rect 149088 614898 149130 615134
rect 149366 614898 149408 615134
rect 149088 614866 149408 614898
rect 179808 615454 180128 615486
rect 179808 615218 179850 615454
rect 180086 615218 180128 615454
rect 179808 615134 180128 615218
rect 179808 614898 179850 615134
rect 180086 614898 180128 615134
rect 179808 614866 180128 614898
rect 210528 615454 210848 615486
rect 210528 615218 210570 615454
rect 210806 615218 210848 615454
rect 210528 615134 210848 615218
rect 210528 614898 210570 615134
rect 210806 614898 210848 615134
rect 210528 614866 210848 614898
rect 241248 615454 241568 615486
rect 241248 615218 241290 615454
rect 241526 615218 241568 615454
rect 241248 615134 241568 615218
rect 241248 614898 241290 615134
rect 241526 614898 241568 615134
rect 241248 614866 241568 614898
rect 271968 615454 272288 615486
rect 271968 615218 272010 615454
rect 272246 615218 272288 615454
rect 271968 615134 272288 615218
rect 271968 614898 272010 615134
rect 272246 614898 272288 615134
rect 271968 614866 272288 614898
rect 302688 615454 303008 615486
rect 302688 615218 302730 615454
rect 302966 615218 303008 615454
rect 302688 615134 303008 615218
rect 302688 614898 302730 615134
rect 302966 614898 303008 615134
rect 302688 614866 303008 614898
rect 333408 615454 333728 615486
rect 333408 615218 333450 615454
rect 333686 615218 333728 615454
rect 333408 615134 333728 615218
rect 333408 614898 333450 615134
rect 333686 614898 333728 615134
rect 333408 614866 333728 614898
rect 364128 615454 364448 615486
rect 364128 615218 364170 615454
rect 364406 615218 364448 615454
rect 364128 615134 364448 615218
rect 364128 614898 364170 615134
rect 364406 614898 364448 615134
rect 364128 614866 364448 614898
rect 394848 615454 395168 615486
rect 394848 615218 394890 615454
rect 395126 615218 395168 615454
rect 394848 615134 395168 615218
rect 394848 614898 394890 615134
rect 395126 614898 395168 615134
rect 394848 614866 395168 614898
rect 425568 615454 425888 615486
rect 425568 615218 425610 615454
rect 425846 615218 425888 615454
rect 425568 615134 425888 615218
rect 425568 614898 425610 615134
rect 425846 614898 425888 615134
rect 425568 614866 425888 614898
rect 456288 615454 456608 615486
rect 456288 615218 456330 615454
rect 456566 615218 456608 615454
rect 456288 615134 456608 615218
rect 456288 614898 456330 615134
rect 456566 614898 456608 615134
rect 456288 614866 456608 614898
rect 487008 615454 487328 615486
rect 487008 615218 487050 615454
rect 487286 615218 487328 615454
rect 487008 615134 487328 615218
rect 487008 614898 487050 615134
rect 487286 614898 487328 615134
rect 487008 614866 487328 614898
rect 517728 615454 518048 615486
rect 517728 615218 517770 615454
rect 518006 615218 518048 615454
rect 517728 615134 518048 615218
rect 517728 614898 517770 615134
rect 518006 614898 518048 615134
rect 517728 614866 518048 614898
rect 548448 615454 548768 615486
rect 548448 615218 548490 615454
rect 548726 615218 548768 615454
rect 548448 615134 548768 615218
rect 548448 614898 548490 615134
rect 548726 614898 548768 615134
rect 548448 614866 548768 614898
rect 24114 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 24734 601774
rect 24114 601454 24734 601538
rect 24114 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 24734 601454
rect 24114 565774 24734 601218
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 41568 583174 41888 583206
rect 41568 582938 41610 583174
rect 41846 582938 41888 583174
rect 41568 582854 41888 582938
rect 41568 582618 41610 582854
rect 41846 582618 41888 582854
rect 41568 582586 41888 582618
rect 72288 583174 72608 583206
rect 72288 582938 72330 583174
rect 72566 582938 72608 583174
rect 72288 582854 72608 582938
rect 72288 582618 72330 582854
rect 72566 582618 72608 582854
rect 72288 582586 72608 582618
rect 103008 583174 103328 583206
rect 103008 582938 103050 583174
rect 103286 582938 103328 583174
rect 103008 582854 103328 582938
rect 103008 582618 103050 582854
rect 103286 582618 103328 582854
rect 103008 582586 103328 582618
rect 133728 583174 134048 583206
rect 133728 582938 133770 583174
rect 134006 582938 134048 583174
rect 133728 582854 134048 582938
rect 133728 582618 133770 582854
rect 134006 582618 134048 582854
rect 133728 582586 134048 582618
rect 164448 583174 164768 583206
rect 164448 582938 164490 583174
rect 164726 582938 164768 583174
rect 164448 582854 164768 582938
rect 164448 582618 164490 582854
rect 164726 582618 164768 582854
rect 164448 582586 164768 582618
rect 195168 583174 195488 583206
rect 195168 582938 195210 583174
rect 195446 582938 195488 583174
rect 195168 582854 195488 582938
rect 195168 582618 195210 582854
rect 195446 582618 195488 582854
rect 195168 582586 195488 582618
rect 225888 583174 226208 583206
rect 225888 582938 225930 583174
rect 226166 582938 226208 583174
rect 225888 582854 226208 582938
rect 225888 582618 225930 582854
rect 226166 582618 226208 582854
rect 225888 582586 226208 582618
rect 256608 583174 256928 583206
rect 256608 582938 256650 583174
rect 256886 582938 256928 583174
rect 256608 582854 256928 582938
rect 256608 582618 256650 582854
rect 256886 582618 256928 582854
rect 256608 582586 256928 582618
rect 287328 583174 287648 583206
rect 287328 582938 287370 583174
rect 287606 582938 287648 583174
rect 287328 582854 287648 582938
rect 287328 582618 287370 582854
rect 287606 582618 287648 582854
rect 287328 582586 287648 582618
rect 318048 583174 318368 583206
rect 318048 582938 318090 583174
rect 318326 582938 318368 583174
rect 318048 582854 318368 582938
rect 318048 582618 318090 582854
rect 318326 582618 318368 582854
rect 318048 582586 318368 582618
rect 348768 583174 349088 583206
rect 348768 582938 348810 583174
rect 349046 582938 349088 583174
rect 348768 582854 349088 582938
rect 348768 582618 348810 582854
rect 349046 582618 349088 582854
rect 348768 582586 349088 582618
rect 379488 583174 379808 583206
rect 379488 582938 379530 583174
rect 379766 582938 379808 583174
rect 379488 582854 379808 582938
rect 379488 582618 379530 582854
rect 379766 582618 379808 582854
rect 379488 582586 379808 582618
rect 410208 583174 410528 583206
rect 410208 582938 410250 583174
rect 410486 582938 410528 583174
rect 410208 582854 410528 582938
rect 410208 582618 410250 582854
rect 410486 582618 410528 582854
rect 410208 582586 410528 582618
rect 440928 583174 441248 583206
rect 440928 582938 440970 583174
rect 441206 582938 441248 583174
rect 440928 582854 441248 582938
rect 440928 582618 440970 582854
rect 441206 582618 441248 582854
rect 440928 582586 441248 582618
rect 471648 583174 471968 583206
rect 471648 582938 471690 583174
rect 471926 582938 471968 583174
rect 471648 582854 471968 582938
rect 471648 582618 471690 582854
rect 471926 582618 471968 582854
rect 471648 582586 471968 582618
rect 502368 583174 502688 583206
rect 502368 582938 502410 583174
rect 502646 582938 502688 583174
rect 502368 582854 502688 582938
rect 502368 582618 502410 582854
rect 502646 582618 502688 582854
rect 502368 582586 502688 582618
rect 533088 583174 533408 583206
rect 533088 582938 533130 583174
rect 533366 582938 533408 583174
rect 533088 582854 533408 582938
rect 533088 582618 533130 582854
rect 533366 582618 533408 582854
rect 533088 582586 533408 582618
rect 26208 579454 26528 579486
rect 26208 579218 26250 579454
rect 26486 579218 26528 579454
rect 26208 579134 26528 579218
rect 26208 578898 26250 579134
rect 26486 578898 26528 579134
rect 26208 578866 26528 578898
rect 56928 579454 57248 579486
rect 56928 579218 56970 579454
rect 57206 579218 57248 579454
rect 56928 579134 57248 579218
rect 56928 578898 56970 579134
rect 57206 578898 57248 579134
rect 56928 578866 57248 578898
rect 87648 579454 87968 579486
rect 87648 579218 87690 579454
rect 87926 579218 87968 579454
rect 87648 579134 87968 579218
rect 87648 578898 87690 579134
rect 87926 578898 87968 579134
rect 87648 578866 87968 578898
rect 118368 579454 118688 579486
rect 118368 579218 118410 579454
rect 118646 579218 118688 579454
rect 118368 579134 118688 579218
rect 118368 578898 118410 579134
rect 118646 578898 118688 579134
rect 118368 578866 118688 578898
rect 149088 579454 149408 579486
rect 149088 579218 149130 579454
rect 149366 579218 149408 579454
rect 149088 579134 149408 579218
rect 149088 578898 149130 579134
rect 149366 578898 149408 579134
rect 149088 578866 149408 578898
rect 179808 579454 180128 579486
rect 179808 579218 179850 579454
rect 180086 579218 180128 579454
rect 179808 579134 180128 579218
rect 179808 578898 179850 579134
rect 180086 578898 180128 579134
rect 179808 578866 180128 578898
rect 210528 579454 210848 579486
rect 210528 579218 210570 579454
rect 210806 579218 210848 579454
rect 210528 579134 210848 579218
rect 210528 578898 210570 579134
rect 210806 578898 210848 579134
rect 210528 578866 210848 578898
rect 241248 579454 241568 579486
rect 241248 579218 241290 579454
rect 241526 579218 241568 579454
rect 241248 579134 241568 579218
rect 241248 578898 241290 579134
rect 241526 578898 241568 579134
rect 241248 578866 241568 578898
rect 271968 579454 272288 579486
rect 271968 579218 272010 579454
rect 272246 579218 272288 579454
rect 271968 579134 272288 579218
rect 271968 578898 272010 579134
rect 272246 578898 272288 579134
rect 271968 578866 272288 578898
rect 302688 579454 303008 579486
rect 302688 579218 302730 579454
rect 302966 579218 303008 579454
rect 302688 579134 303008 579218
rect 302688 578898 302730 579134
rect 302966 578898 303008 579134
rect 302688 578866 303008 578898
rect 333408 579454 333728 579486
rect 333408 579218 333450 579454
rect 333686 579218 333728 579454
rect 333408 579134 333728 579218
rect 333408 578898 333450 579134
rect 333686 578898 333728 579134
rect 333408 578866 333728 578898
rect 364128 579454 364448 579486
rect 364128 579218 364170 579454
rect 364406 579218 364448 579454
rect 364128 579134 364448 579218
rect 364128 578898 364170 579134
rect 364406 578898 364448 579134
rect 364128 578866 364448 578898
rect 394848 579454 395168 579486
rect 394848 579218 394890 579454
rect 395126 579218 395168 579454
rect 394848 579134 395168 579218
rect 394848 578898 394890 579134
rect 395126 578898 395168 579134
rect 394848 578866 395168 578898
rect 425568 579454 425888 579486
rect 425568 579218 425610 579454
rect 425846 579218 425888 579454
rect 425568 579134 425888 579218
rect 425568 578898 425610 579134
rect 425846 578898 425888 579134
rect 425568 578866 425888 578898
rect 456288 579454 456608 579486
rect 456288 579218 456330 579454
rect 456566 579218 456608 579454
rect 456288 579134 456608 579218
rect 456288 578898 456330 579134
rect 456566 578898 456608 579134
rect 456288 578866 456608 578898
rect 487008 579454 487328 579486
rect 487008 579218 487050 579454
rect 487286 579218 487328 579454
rect 487008 579134 487328 579218
rect 487008 578898 487050 579134
rect 487286 578898 487328 579134
rect 487008 578866 487328 578898
rect 517728 579454 518048 579486
rect 517728 579218 517770 579454
rect 518006 579218 518048 579454
rect 517728 579134 518048 579218
rect 517728 578898 517770 579134
rect 518006 578898 518048 579134
rect 517728 578866 518048 578898
rect 548448 579454 548768 579486
rect 548448 579218 548490 579454
rect 548726 579218 548768 579454
rect 548448 579134 548768 579218
rect 548448 578898 548490 579134
rect 548726 578898 548768 579134
rect 548448 578866 548768 578898
rect 24114 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 24734 565774
rect 24114 565454 24734 565538
rect 24114 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 24734 565454
rect 24114 529774 24734 565218
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 41568 547174 41888 547206
rect 41568 546938 41610 547174
rect 41846 546938 41888 547174
rect 41568 546854 41888 546938
rect 41568 546618 41610 546854
rect 41846 546618 41888 546854
rect 41568 546586 41888 546618
rect 72288 547174 72608 547206
rect 72288 546938 72330 547174
rect 72566 546938 72608 547174
rect 72288 546854 72608 546938
rect 72288 546618 72330 546854
rect 72566 546618 72608 546854
rect 72288 546586 72608 546618
rect 103008 547174 103328 547206
rect 103008 546938 103050 547174
rect 103286 546938 103328 547174
rect 103008 546854 103328 546938
rect 103008 546618 103050 546854
rect 103286 546618 103328 546854
rect 103008 546586 103328 546618
rect 133728 547174 134048 547206
rect 133728 546938 133770 547174
rect 134006 546938 134048 547174
rect 133728 546854 134048 546938
rect 133728 546618 133770 546854
rect 134006 546618 134048 546854
rect 133728 546586 134048 546618
rect 164448 547174 164768 547206
rect 164448 546938 164490 547174
rect 164726 546938 164768 547174
rect 164448 546854 164768 546938
rect 164448 546618 164490 546854
rect 164726 546618 164768 546854
rect 164448 546586 164768 546618
rect 195168 547174 195488 547206
rect 195168 546938 195210 547174
rect 195446 546938 195488 547174
rect 195168 546854 195488 546938
rect 195168 546618 195210 546854
rect 195446 546618 195488 546854
rect 195168 546586 195488 546618
rect 225888 547174 226208 547206
rect 225888 546938 225930 547174
rect 226166 546938 226208 547174
rect 225888 546854 226208 546938
rect 225888 546618 225930 546854
rect 226166 546618 226208 546854
rect 225888 546586 226208 546618
rect 256608 547174 256928 547206
rect 256608 546938 256650 547174
rect 256886 546938 256928 547174
rect 256608 546854 256928 546938
rect 256608 546618 256650 546854
rect 256886 546618 256928 546854
rect 256608 546586 256928 546618
rect 287328 547174 287648 547206
rect 287328 546938 287370 547174
rect 287606 546938 287648 547174
rect 287328 546854 287648 546938
rect 287328 546618 287370 546854
rect 287606 546618 287648 546854
rect 287328 546586 287648 546618
rect 318048 547174 318368 547206
rect 318048 546938 318090 547174
rect 318326 546938 318368 547174
rect 318048 546854 318368 546938
rect 318048 546618 318090 546854
rect 318326 546618 318368 546854
rect 318048 546586 318368 546618
rect 348768 547174 349088 547206
rect 348768 546938 348810 547174
rect 349046 546938 349088 547174
rect 348768 546854 349088 546938
rect 348768 546618 348810 546854
rect 349046 546618 349088 546854
rect 348768 546586 349088 546618
rect 379488 547174 379808 547206
rect 379488 546938 379530 547174
rect 379766 546938 379808 547174
rect 379488 546854 379808 546938
rect 379488 546618 379530 546854
rect 379766 546618 379808 546854
rect 379488 546586 379808 546618
rect 410208 547174 410528 547206
rect 410208 546938 410250 547174
rect 410486 546938 410528 547174
rect 410208 546854 410528 546938
rect 410208 546618 410250 546854
rect 410486 546618 410528 546854
rect 410208 546586 410528 546618
rect 440928 547174 441248 547206
rect 440928 546938 440970 547174
rect 441206 546938 441248 547174
rect 440928 546854 441248 546938
rect 440928 546618 440970 546854
rect 441206 546618 441248 546854
rect 440928 546586 441248 546618
rect 471648 547174 471968 547206
rect 471648 546938 471690 547174
rect 471926 546938 471968 547174
rect 471648 546854 471968 546938
rect 471648 546618 471690 546854
rect 471926 546618 471968 546854
rect 471648 546586 471968 546618
rect 502368 547174 502688 547206
rect 502368 546938 502410 547174
rect 502646 546938 502688 547174
rect 502368 546854 502688 546938
rect 502368 546618 502410 546854
rect 502646 546618 502688 546854
rect 502368 546586 502688 546618
rect 533088 547174 533408 547206
rect 533088 546938 533130 547174
rect 533366 546938 533408 547174
rect 533088 546854 533408 546938
rect 533088 546618 533130 546854
rect 533366 546618 533408 546854
rect 533088 546586 533408 546618
rect 26208 543454 26528 543486
rect 26208 543218 26250 543454
rect 26486 543218 26528 543454
rect 26208 543134 26528 543218
rect 26208 542898 26250 543134
rect 26486 542898 26528 543134
rect 26208 542866 26528 542898
rect 56928 543454 57248 543486
rect 56928 543218 56970 543454
rect 57206 543218 57248 543454
rect 56928 543134 57248 543218
rect 56928 542898 56970 543134
rect 57206 542898 57248 543134
rect 56928 542866 57248 542898
rect 87648 543454 87968 543486
rect 87648 543218 87690 543454
rect 87926 543218 87968 543454
rect 87648 543134 87968 543218
rect 87648 542898 87690 543134
rect 87926 542898 87968 543134
rect 87648 542866 87968 542898
rect 118368 543454 118688 543486
rect 118368 543218 118410 543454
rect 118646 543218 118688 543454
rect 118368 543134 118688 543218
rect 118368 542898 118410 543134
rect 118646 542898 118688 543134
rect 118368 542866 118688 542898
rect 149088 543454 149408 543486
rect 149088 543218 149130 543454
rect 149366 543218 149408 543454
rect 149088 543134 149408 543218
rect 149088 542898 149130 543134
rect 149366 542898 149408 543134
rect 149088 542866 149408 542898
rect 179808 543454 180128 543486
rect 179808 543218 179850 543454
rect 180086 543218 180128 543454
rect 179808 543134 180128 543218
rect 179808 542898 179850 543134
rect 180086 542898 180128 543134
rect 179808 542866 180128 542898
rect 210528 543454 210848 543486
rect 210528 543218 210570 543454
rect 210806 543218 210848 543454
rect 210528 543134 210848 543218
rect 210528 542898 210570 543134
rect 210806 542898 210848 543134
rect 210528 542866 210848 542898
rect 241248 543454 241568 543486
rect 241248 543218 241290 543454
rect 241526 543218 241568 543454
rect 241248 543134 241568 543218
rect 241248 542898 241290 543134
rect 241526 542898 241568 543134
rect 241248 542866 241568 542898
rect 271968 543454 272288 543486
rect 271968 543218 272010 543454
rect 272246 543218 272288 543454
rect 271968 543134 272288 543218
rect 271968 542898 272010 543134
rect 272246 542898 272288 543134
rect 271968 542866 272288 542898
rect 302688 543454 303008 543486
rect 302688 543218 302730 543454
rect 302966 543218 303008 543454
rect 302688 543134 303008 543218
rect 302688 542898 302730 543134
rect 302966 542898 303008 543134
rect 302688 542866 303008 542898
rect 333408 543454 333728 543486
rect 333408 543218 333450 543454
rect 333686 543218 333728 543454
rect 333408 543134 333728 543218
rect 333408 542898 333450 543134
rect 333686 542898 333728 543134
rect 333408 542866 333728 542898
rect 364128 543454 364448 543486
rect 364128 543218 364170 543454
rect 364406 543218 364448 543454
rect 364128 543134 364448 543218
rect 364128 542898 364170 543134
rect 364406 542898 364448 543134
rect 364128 542866 364448 542898
rect 394848 543454 395168 543486
rect 394848 543218 394890 543454
rect 395126 543218 395168 543454
rect 394848 543134 395168 543218
rect 394848 542898 394890 543134
rect 395126 542898 395168 543134
rect 394848 542866 395168 542898
rect 425568 543454 425888 543486
rect 425568 543218 425610 543454
rect 425846 543218 425888 543454
rect 425568 543134 425888 543218
rect 425568 542898 425610 543134
rect 425846 542898 425888 543134
rect 425568 542866 425888 542898
rect 456288 543454 456608 543486
rect 456288 543218 456330 543454
rect 456566 543218 456608 543454
rect 456288 543134 456608 543218
rect 456288 542898 456330 543134
rect 456566 542898 456608 543134
rect 456288 542866 456608 542898
rect 487008 543454 487328 543486
rect 487008 543218 487050 543454
rect 487286 543218 487328 543454
rect 487008 543134 487328 543218
rect 487008 542898 487050 543134
rect 487286 542898 487328 543134
rect 487008 542866 487328 542898
rect 517728 543454 518048 543486
rect 517728 543218 517770 543454
rect 518006 543218 518048 543454
rect 517728 543134 518048 543218
rect 517728 542898 517770 543134
rect 518006 542898 518048 543134
rect 517728 542866 518048 542898
rect 548448 543454 548768 543486
rect 548448 543218 548490 543454
rect 548726 543218 548768 543454
rect 548448 543134 548768 543218
rect 548448 542898 548490 543134
rect 548726 542898 548768 543134
rect 548448 542866 548768 542898
rect 24114 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 24734 529774
rect 24114 529454 24734 529538
rect 24114 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 24734 529454
rect 24114 493774 24734 529218
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 41568 511174 41888 511206
rect 41568 510938 41610 511174
rect 41846 510938 41888 511174
rect 41568 510854 41888 510938
rect 41568 510618 41610 510854
rect 41846 510618 41888 510854
rect 41568 510586 41888 510618
rect 72288 511174 72608 511206
rect 72288 510938 72330 511174
rect 72566 510938 72608 511174
rect 72288 510854 72608 510938
rect 72288 510618 72330 510854
rect 72566 510618 72608 510854
rect 72288 510586 72608 510618
rect 103008 511174 103328 511206
rect 103008 510938 103050 511174
rect 103286 510938 103328 511174
rect 103008 510854 103328 510938
rect 103008 510618 103050 510854
rect 103286 510618 103328 510854
rect 103008 510586 103328 510618
rect 133728 511174 134048 511206
rect 133728 510938 133770 511174
rect 134006 510938 134048 511174
rect 133728 510854 134048 510938
rect 133728 510618 133770 510854
rect 134006 510618 134048 510854
rect 133728 510586 134048 510618
rect 164448 511174 164768 511206
rect 164448 510938 164490 511174
rect 164726 510938 164768 511174
rect 164448 510854 164768 510938
rect 164448 510618 164490 510854
rect 164726 510618 164768 510854
rect 164448 510586 164768 510618
rect 195168 511174 195488 511206
rect 195168 510938 195210 511174
rect 195446 510938 195488 511174
rect 195168 510854 195488 510938
rect 195168 510618 195210 510854
rect 195446 510618 195488 510854
rect 195168 510586 195488 510618
rect 225888 511174 226208 511206
rect 225888 510938 225930 511174
rect 226166 510938 226208 511174
rect 225888 510854 226208 510938
rect 225888 510618 225930 510854
rect 226166 510618 226208 510854
rect 225888 510586 226208 510618
rect 256608 511174 256928 511206
rect 256608 510938 256650 511174
rect 256886 510938 256928 511174
rect 256608 510854 256928 510938
rect 256608 510618 256650 510854
rect 256886 510618 256928 510854
rect 256608 510586 256928 510618
rect 287328 511174 287648 511206
rect 287328 510938 287370 511174
rect 287606 510938 287648 511174
rect 287328 510854 287648 510938
rect 287328 510618 287370 510854
rect 287606 510618 287648 510854
rect 287328 510586 287648 510618
rect 318048 511174 318368 511206
rect 318048 510938 318090 511174
rect 318326 510938 318368 511174
rect 318048 510854 318368 510938
rect 318048 510618 318090 510854
rect 318326 510618 318368 510854
rect 318048 510586 318368 510618
rect 348768 511174 349088 511206
rect 348768 510938 348810 511174
rect 349046 510938 349088 511174
rect 348768 510854 349088 510938
rect 348768 510618 348810 510854
rect 349046 510618 349088 510854
rect 348768 510586 349088 510618
rect 379488 511174 379808 511206
rect 379488 510938 379530 511174
rect 379766 510938 379808 511174
rect 379488 510854 379808 510938
rect 379488 510618 379530 510854
rect 379766 510618 379808 510854
rect 379488 510586 379808 510618
rect 410208 511174 410528 511206
rect 410208 510938 410250 511174
rect 410486 510938 410528 511174
rect 410208 510854 410528 510938
rect 410208 510618 410250 510854
rect 410486 510618 410528 510854
rect 410208 510586 410528 510618
rect 440928 511174 441248 511206
rect 440928 510938 440970 511174
rect 441206 510938 441248 511174
rect 440928 510854 441248 510938
rect 440928 510618 440970 510854
rect 441206 510618 441248 510854
rect 440928 510586 441248 510618
rect 471648 511174 471968 511206
rect 471648 510938 471690 511174
rect 471926 510938 471968 511174
rect 471648 510854 471968 510938
rect 471648 510618 471690 510854
rect 471926 510618 471968 510854
rect 471648 510586 471968 510618
rect 502368 511174 502688 511206
rect 502368 510938 502410 511174
rect 502646 510938 502688 511174
rect 502368 510854 502688 510938
rect 502368 510618 502410 510854
rect 502646 510618 502688 510854
rect 502368 510586 502688 510618
rect 533088 511174 533408 511206
rect 533088 510938 533130 511174
rect 533366 510938 533408 511174
rect 533088 510854 533408 510938
rect 533088 510618 533130 510854
rect 533366 510618 533408 510854
rect 533088 510586 533408 510618
rect 26208 507454 26528 507486
rect 26208 507218 26250 507454
rect 26486 507218 26528 507454
rect 26208 507134 26528 507218
rect 26208 506898 26250 507134
rect 26486 506898 26528 507134
rect 26208 506866 26528 506898
rect 56928 507454 57248 507486
rect 56928 507218 56970 507454
rect 57206 507218 57248 507454
rect 56928 507134 57248 507218
rect 56928 506898 56970 507134
rect 57206 506898 57248 507134
rect 56928 506866 57248 506898
rect 87648 507454 87968 507486
rect 87648 507218 87690 507454
rect 87926 507218 87968 507454
rect 87648 507134 87968 507218
rect 87648 506898 87690 507134
rect 87926 506898 87968 507134
rect 87648 506866 87968 506898
rect 118368 507454 118688 507486
rect 118368 507218 118410 507454
rect 118646 507218 118688 507454
rect 118368 507134 118688 507218
rect 118368 506898 118410 507134
rect 118646 506898 118688 507134
rect 118368 506866 118688 506898
rect 149088 507454 149408 507486
rect 149088 507218 149130 507454
rect 149366 507218 149408 507454
rect 149088 507134 149408 507218
rect 149088 506898 149130 507134
rect 149366 506898 149408 507134
rect 149088 506866 149408 506898
rect 179808 507454 180128 507486
rect 179808 507218 179850 507454
rect 180086 507218 180128 507454
rect 179808 507134 180128 507218
rect 179808 506898 179850 507134
rect 180086 506898 180128 507134
rect 179808 506866 180128 506898
rect 210528 507454 210848 507486
rect 210528 507218 210570 507454
rect 210806 507218 210848 507454
rect 210528 507134 210848 507218
rect 210528 506898 210570 507134
rect 210806 506898 210848 507134
rect 210528 506866 210848 506898
rect 241248 507454 241568 507486
rect 241248 507218 241290 507454
rect 241526 507218 241568 507454
rect 241248 507134 241568 507218
rect 241248 506898 241290 507134
rect 241526 506898 241568 507134
rect 241248 506866 241568 506898
rect 271968 507454 272288 507486
rect 271968 507218 272010 507454
rect 272246 507218 272288 507454
rect 271968 507134 272288 507218
rect 271968 506898 272010 507134
rect 272246 506898 272288 507134
rect 271968 506866 272288 506898
rect 302688 507454 303008 507486
rect 302688 507218 302730 507454
rect 302966 507218 303008 507454
rect 302688 507134 303008 507218
rect 302688 506898 302730 507134
rect 302966 506898 303008 507134
rect 302688 506866 303008 506898
rect 333408 507454 333728 507486
rect 333408 507218 333450 507454
rect 333686 507218 333728 507454
rect 333408 507134 333728 507218
rect 333408 506898 333450 507134
rect 333686 506898 333728 507134
rect 333408 506866 333728 506898
rect 364128 507454 364448 507486
rect 364128 507218 364170 507454
rect 364406 507218 364448 507454
rect 364128 507134 364448 507218
rect 364128 506898 364170 507134
rect 364406 506898 364448 507134
rect 364128 506866 364448 506898
rect 394848 507454 395168 507486
rect 394848 507218 394890 507454
rect 395126 507218 395168 507454
rect 394848 507134 395168 507218
rect 394848 506898 394890 507134
rect 395126 506898 395168 507134
rect 394848 506866 395168 506898
rect 425568 507454 425888 507486
rect 425568 507218 425610 507454
rect 425846 507218 425888 507454
rect 425568 507134 425888 507218
rect 425568 506898 425610 507134
rect 425846 506898 425888 507134
rect 425568 506866 425888 506898
rect 456288 507454 456608 507486
rect 456288 507218 456330 507454
rect 456566 507218 456608 507454
rect 456288 507134 456608 507218
rect 456288 506898 456330 507134
rect 456566 506898 456608 507134
rect 456288 506866 456608 506898
rect 487008 507454 487328 507486
rect 487008 507218 487050 507454
rect 487286 507218 487328 507454
rect 487008 507134 487328 507218
rect 487008 506898 487050 507134
rect 487286 506898 487328 507134
rect 487008 506866 487328 506898
rect 517728 507454 518048 507486
rect 517728 507218 517770 507454
rect 518006 507218 518048 507454
rect 517728 507134 518048 507218
rect 517728 506898 517770 507134
rect 518006 506898 518048 507134
rect 517728 506866 518048 506898
rect 548448 507454 548768 507486
rect 548448 507218 548490 507454
rect 548726 507218 548768 507454
rect 548448 507134 548768 507218
rect 548448 506898 548490 507134
rect 548726 506898 548768 507134
rect 548448 506866 548768 506898
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 41568 475174 41888 475206
rect 41568 474938 41610 475174
rect 41846 474938 41888 475174
rect 41568 474854 41888 474938
rect 41568 474618 41610 474854
rect 41846 474618 41888 474854
rect 41568 474586 41888 474618
rect 72288 475174 72608 475206
rect 72288 474938 72330 475174
rect 72566 474938 72608 475174
rect 72288 474854 72608 474938
rect 72288 474618 72330 474854
rect 72566 474618 72608 474854
rect 72288 474586 72608 474618
rect 103008 475174 103328 475206
rect 103008 474938 103050 475174
rect 103286 474938 103328 475174
rect 103008 474854 103328 474938
rect 103008 474618 103050 474854
rect 103286 474618 103328 474854
rect 103008 474586 103328 474618
rect 133728 475174 134048 475206
rect 133728 474938 133770 475174
rect 134006 474938 134048 475174
rect 133728 474854 134048 474938
rect 133728 474618 133770 474854
rect 134006 474618 134048 474854
rect 133728 474586 134048 474618
rect 164448 475174 164768 475206
rect 164448 474938 164490 475174
rect 164726 474938 164768 475174
rect 164448 474854 164768 474938
rect 164448 474618 164490 474854
rect 164726 474618 164768 474854
rect 164448 474586 164768 474618
rect 195168 475174 195488 475206
rect 195168 474938 195210 475174
rect 195446 474938 195488 475174
rect 195168 474854 195488 474938
rect 195168 474618 195210 474854
rect 195446 474618 195488 474854
rect 195168 474586 195488 474618
rect 225888 475174 226208 475206
rect 225888 474938 225930 475174
rect 226166 474938 226208 475174
rect 225888 474854 226208 474938
rect 225888 474618 225930 474854
rect 226166 474618 226208 474854
rect 225888 474586 226208 474618
rect 256608 475174 256928 475206
rect 256608 474938 256650 475174
rect 256886 474938 256928 475174
rect 256608 474854 256928 474938
rect 256608 474618 256650 474854
rect 256886 474618 256928 474854
rect 256608 474586 256928 474618
rect 287328 475174 287648 475206
rect 287328 474938 287370 475174
rect 287606 474938 287648 475174
rect 287328 474854 287648 474938
rect 287328 474618 287370 474854
rect 287606 474618 287648 474854
rect 287328 474586 287648 474618
rect 318048 475174 318368 475206
rect 318048 474938 318090 475174
rect 318326 474938 318368 475174
rect 318048 474854 318368 474938
rect 318048 474618 318090 474854
rect 318326 474618 318368 474854
rect 318048 474586 318368 474618
rect 348768 475174 349088 475206
rect 348768 474938 348810 475174
rect 349046 474938 349088 475174
rect 348768 474854 349088 474938
rect 348768 474618 348810 474854
rect 349046 474618 349088 474854
rect 348768 474586 349088 474618
rect 379488 475174 379808 475206
rect 379488 474938 379530 475174
rect 379766 474938 379808 475174
rect 379488 474854 379808 474938
rect 379488 474618 379530 474854
rect 379766 474618 379808 474854
rect 379488 474586 379808 474618
rect 410208 475174 410528 475206
rect 410208 474938 410250 475174
rect 410486 474938 410528 475174
rect 410208 474854 410528 474938
rect 410208 474618 410250 474854
rect 410486 474618 410528 474854
rect 410208 474586 410528 474618
rect 440928 475174 441248 475206
rect 440928 474938 440970 475174
rect 441206 474938 441248 475174
rect 440928 474854 441248 474938
rect 440928 474618 440970 474854
rect 441206 474618 441248 474854
rect 440928 474586 441248 474618
rect 471648 475174 471968 475206
rect 471648 474938 471690 475174
rect 471926 474938 471968 475174
rect 471648 474854 471968 474938
rect 471648 474618 471690 474854
rect 471926 474618 471968 474854
rect 471648 474586 471968 474618
rect 502368 475174 502688 475206
rect 502368 474938 502410 475174
rect 502646 474938 502688 475174
rect 502368 474854 502688 474938
rect 502368 474618 502410 474854
rect 502646 474618 502688 474854
rect 502368 474586 502688 474618
rect 533088 475174 533408 475206
rect 533088 474938 533130 475174
rect 533366 474938 533408 475174
rect 533088 474854 533408 474938
rect 533088 474618 533130 474854
rect 533366 474618 533408 474854
rect 533088 474586 533408 474618
rect 26208 471454 26528 471486
rect 26208 471218 26250 471454
rect 26486 471218 26528 471454
rect 26208 471134 26528 471218
rect 26208 470898 26250 471134
rect 26486 470898 26528 471134
rect 26208 470866 26528 470898
rect 56928 471454 57248 471486
rect 56928 471218 56970 471454
rect 57206 471218 57248 471454
rect 56928 471134 57248 471218
rect 56928 470898 56970 471134
rect 57206 470898 57248 471134
rect 56928 470866 57248 470898
rect 87648 471454 87968 471486
rect 87648 471218 87690 471454
rect 87926 471218 87968 471454
rect 87648 471134 87968 471218
rect 87648 470898 87690 471134
rect 87926 470898 87968 471134
rect 87648 470866 87968 470898
rect 118368 471454 118688 471486
rect 118368 471218 118410 471454
rect 118646 471218 118688 471454
rect 118368 471134 118688 471218
rect 118368 470898 118410 471134
rect 118646 470898 118688 471134
rect 118368 470866 118688 470898
rect 149088 471454 149408 471486
rect 149088 471218 149130 471454
rect 149366 471218 149408 471454
rect 149088 471134 149408 471218
rect 149088 470898 149130 471134
rect 149366 470898 149408 471134
rect 149088 470866 149408 470898
rect 179808 471454 180128 471486
rect 179808 471218 179850 471454
rect 180086 471218 180128 471454
rect 179808 471134 180128 471218
rect 179808 470898 179850 471134
rect 180086 470898 180128 471134
rect 179808 470866 180128 470898
rect 210528 471454 210848 471486
rect 210528 471218 210570 471454
rect 210806 471218 210848 471454
rect 210528 471134 210848 471218
rect 210528 470898 210570 471134
rect 210806 470898 210848 471134
rect 210528 470866 210848 470898
rect 241248 471454 241568 471486
rect 241248 471218 241290 471454
rect 241526 471218 241568 471454
rect 241248 471134 241568 471218
rect 241248 470898 241290 471134
rect 241526 470898 241568 471134
rect 241248 470866 241568 470898
rect 271968 471454 272288 471486
rect 271968 471218 272010 471454
rect 272246 471218 272288 471454
rect 271968 471134 272288 471218
rect 271968 470898 272010 471134
rect 272246 470898 272288 471134
rect 271968 470866 272288 470898
rect 302688 471454 303008 471486
rect 302688 471218 302730 471454
rect 302966 471218 303008 471454
rect 302688 471134 303008 471218
rect 302688 470898 302730 471134
rect 302966 470898 303008 471134
rect 302688 470866 303008 470898
rect 333408 471454 333728 471486
rect 333408 471218 333450 471454
rect 333686 471218 333728 471454
rect 333408 471134 333728 471218
rect 333408 470898 333450 471134
rect 333686 470898 333728 471134
rect 333408 470866 333728 470898
rect 364128 471454 364448 471486
rect 364128 471218 364170 471454
rect 364406 471218 364448 471454
rect 364128 471134 364448 471218
rect 364128 470898 364170 471134
rect 364406 470898 364448 471134
rect 364128 470866 364448 470898
rect 394848 471454 395168 471486
rect 394848 471218 394890 471454
rect 395126 471218 395168 471454
rect 394848 471134 395168 471218
rect 394848 470898 394890 471134
rect 395126 470898 395168 471134
rect 394848 470866 395168 470898
rect 425568 471454 425888 471486
rect 425568 471218 425610 471454
rect 425846 471218 425888 471454
rect 425568 471134 425888 471218
rect 425568 470898 425610 471134
rect 425846 470898 425888 471134
rect 425568 470866 425888 470898
rect 456288 471454 456608 471486
rect 456288 471218 456330 471454
rect 456566 471218 456608 471454
rect 456288 471134 456608 471218
rect 456288 470898 456330 471134
rect 456566 470898 456608 471134
rect 456288 470866 456608 470898
rect 487008 471454 487328 471486
rect 487008 471218 487050 471454
rect 487286 471218 487328 471454
rect 487008 471134 487328 471218
rect 487008 470898 487050 471134
rect 487286 470898 487328 471134
rect 487008 470866 487328 470898
rect 517728 471454 518048 471486
rect 517728 471218 517770 471454
rect 518006 471218 518048 471454
rect 517728 471134 518048 471218
rect 517728 470898 517770 471134
rect 518006 470898 518048 471134
rect 517728 470866 518048 470898
rect 548448 471454 548768 471486
rect 548448 471218 548490 471454
rect 548726 471218 548768 471454
rect 548448 471134 548768 471218
rect 548448 470898 548490 471134
rect 548726 470898 548768 471134
rect 548448 470866 548768 470898
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 421774 24734 457218
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 41568 439174 41888 439206
rect 41568 438938 41610 439174
rect 41846 438938 41888 439174
rect 41568 438854 41888 438938
rect 41568 438618 41610 438854
rect 41846 438618 41888 438854
rect 41568 438586 41888 438618
rect 72288 439174 72608 439206
rect 72288 438938 72330 439174
rect 72566 438938 72608 439174
rect 72288 438854 72608 438938
rect 72288 438618 72330 438854
rect 72566 438618 72608 438854
rect 72288 438586 72608 438618
rect 103008 439174 103328 439206
rect 103008 438938 103050 439174
rect 103286 438938 103328 439174
rect 103008 438854 103328 438938
rect 103008 438618 103050 438854
rect 103286 438618 103328 438854
rect 103008 438586 103328 438618
rect 133728 439174 134048 439206
rect 133728 438938 133770 439174
rect 134006 438938 134048 439174
rect 133728 438854 134048 438938
rect 133728 438618 133770 438854
rect 134006 438618 134048 438854
rect 133728 438586 134048 438618
rect 164448 439174 164768 439206
rect 164448 438938 164490 439174
rect 164726 438938 164768 439174
rect 164448 438854 164768 438938
rect 164448 438618 164490 438854
rect 164726 438618 164768 438854
rect 164448 438586 164768 438618
rect 195168 439174 195488 439206
rect 195168 438938 195210 439174
rect 195446 438938 195488 439174
rect 195168 438854 195488 438938
rect 195168 438618 195210 438854
rect 195446 438618 195488 438854
rect 195168 438586 195488 438618
rect 225888 439174 226208 439206
rect 225888 438938 225930 439174
rect 226166 438938 226208 439174
rect 225888 438854 226208 438938
rect 225888 438618 225930 438854
rect 226166 438618 226208 438854
rect 225888 438586 226208 438618
rect 256608 439174 256928 439206
rect 256608 438938 256650 439174
rect 256886 438938 256928 439174
rect 256608 438854 256928 438938
rect 256608 438618 256650 438854
rect 256886 438618 256928 438854
rect 256608 438586 256928 438618
rect 287328 439174 287648 439206
rect 287328 438938 287370 439174
rect 287606 438938 287648 439174
rect 287328 438854 287648 438938
rect 287328 438618 287370 438854
rect 287606 438618 287648 438854
rect 287328 438586 287648 438618
rect 318048 439174 318368 439206
rect 318048 438938 318090 439174
rect 318326 438938 318368 439174
rect 318048 438854 318368 438938
rect 318048 438618 318090 438854
rect 318326 438618 318368 438854
rect 318048 438586 318368 438618
rect 348768 439174 349088 439206
rect 348768 438938 348810 439174
rect 349046 438938 349088 439174
rect 348768 438854 349088 438938
rect 348768 438618 348810 438854
rect 349046 438618 349088 438854
rect 348768 438586 349088 438618
rect 379488 439174 379808 439206
rect 379488 438938 379530 439174
rect 379766 438938 379808 439174
rect 379488 438854 379808 438938
rect 379488 438618 379530 438854
rect 379766 438618 379808 438854
rect 379488 438586 379808 438618
rect 410208 439174 410528 439206
rect 410208 438938 410250 439174
rect 410486 438938 410528 439174
rect 410208 438854 410528 438938
rect 410208 438618 410250 438854
rect 410486 438618 410528 438854
rect 410208 438586 410528 438618
rect 440928 439174 441248 439206
rect 440928 438938 440970 439174
rect 441206 438938 441248 439174
rect 440928 438854 441248 438938
rect 440928 438618 440970 438854
rect 441206 438618 441248 438854
rect 440928 438586 441248 438618
rect 471648 439174 471968 439206
rect 471648 438938 471690 439174
rect 471926 438938 471968 439174
rect 471648 438854 471968 438938
rect 471648 438618 471690 438854
rect 471926 438618 471968 438854
rect 471648 438586 471968 438618
rect 502368 439174 502688 439206
rect 502368 438938 502410 439174
rect 502646 438938 502688 439174
rect 502368 438854 502688 438938
rect 502368 438618 502410 438854
rect 502646 438618 502688 438854
rect 502368 438586 502688 438618
rect 533088 439174 533408 439206
rect 533088 438938 533130 439174
rect 533366 438938 533408 439174
rect 533088 438854 533408 438938
rect 533088 438618 533130 438854
rect 533366 438618 533408 438854
rect 533088 438586 533408 438618
rect 26208 435454 26528 435486
rect 26208 435218 26250 435454
rect 26486 435218 26528 435454
rect 26208 435134 26528 435218
rect 26208 434898 26250 435134
rect 26486 434898 26528 435134
rect 26208 434866 26528 434898
rect 56928 435454 57248 435486
rect 56928 435218 56970 435454
rect 57206 435218 57248 435454
rect 56928 435134 57248 435218
rect 56928 434898 56970 435134
rect 57206 434898 57248 435134
rect 56928 434866 57248 434898
rect 87648 435454 87968 435486
rect 87648 435218 87690 435454
rect 87926 435218 87968 435454
rect 87648 435134 87968 435218
rect 87648 434898 87690 435134
rect 87926 434898 87968 435134
rect 87648 434866 87968 434898
rect 118368 435454 118688 435486
rect 118368 435218 118410 435454
rect 118646 435218 118688 435454
rect 118368 435134 118688 435218
rect 118368 434898 118410 435134
rect 118646 434898 118688 435134
rect 118368 434866 118688 434898
rect 149088 435454 149408 435486
rect 149088 435218 149130 435454
rect 149366 435218 149408 435454
rect 149088 435134 149408 435218
rect 149088 434898 149130 435134
rect 149366 434898 149408 435134
rect 149088 434866 149408 434898
rect 179808 435454 180128 435486
rect 179808 435218 179850 435454
rect 180086 435218 180128 435454
rect 179808 435134 180128 435218
rect 179808 434898 179850 435134
rect 180086 434898 180128 435134
rect 179808 434866 180128 434898
rect 210528 435454 210848 435486
rect 210528 435218 210570 435454
rect 210806 435218 210848 435454
rect 210528 435134 210848 435218
rect 210528 434898 210570 435134
rect 210806 434898 210848 435134
rect 210528 434866 210848 434898
rect 241248 435454 241568 435486
rect 241248 435218 241290 435454
rect 241526 435218 241568 435454
rect 241248 435134 241568 435218
rect 241248 434898 241290 435134
rect 241526 434898 241568 435134
rect 241248 434866 241568 434898
rect 271968 435454 272288 435486
rect 271968 435218 272010 435454
rect 272246 435218 272288 435454
rect 271968 435134 272288 435218
rect 271968 434898 272010 435134
rect 272246 434898 272288 435134
rect 271968 434866 272288 434898
rect 302688 435454 303008 435486
rect 302688 435218 302730 435454
rect 302966 435218 303008 435454
rect 302688 435134 303008 435218
rect 302688 434898 302730 435134
rect 302966 434898 303008 435134
rect 302688 434866 303008 434898
rect 333408 435454 333728 435486
rect 333408 435218 333450 435454
rect 333686 435218 333728 435454
rect 333408 435134 333728 435218
rect 333408 434898 333450 435134
rect 333686 434898 333728 435134
rect 333408 434866 333728 434898
rect 364128 435454 364448 435486
rect 364128 435218 364170 435454
rect 364406 435218 364448 435454
rect 364128 435134 364448 435218
rect 364128 434898 364170 435134
rect 364406 434898 364448 435134
rect 364128 434866 364448 434898
rect 394848 435454 395168 435486
rect 394848 435218 394890 435454
rect 395126 435218 395168 435454
rect 394848 435134 395168 435218
rect 394848 434898 394890 435134
rect 395126 434898 395168 435134
rect 394848 434866 395168 434898
rect 425568 435454 425888 435486
rect 425568 435218 425610 435454
rect 425846 435218 425888 435454
rect 425568 435134 425888 435218
rect 425568 434898 425610 435134
rect 425846 434898 425888 435134
rect 425568 434866 425888 434898
rect 456288 435454 456608 435486
rect 456288 435218 456330 435454
rect 456566 435218 456608 435454
rect 456288 435134 456608 435218
rect 456288 434898 456330 435134
rect 456566 434898 456608 435134
rect 456288 434866 456608 434898
rect 487008 435454 487328 435486
rect 487008 435218 487050 435454
rect 487286 435218 487328 435454
rect 487008 435134 487328 435218
rect 487008 434898 487050 435134
rect 487286 434898 487328 435134
rect 487008 434866 487328 434898
rect 517728 435454 518048 435486
rect 517728 435218 517770 435454
rect 518006 435218 518048 435454
rect 517728 435134 518048 435218
rect 517728 434898 517770 435134
rect 518006 434898 518048 435134
rect 517728 434866 518048 434898
rect 548448 435454 548768 435486
rect 548448 435218 548490 435454
rect 548726 435218 548768 435454
rect 548448 435134 548768 435218
rect 548448 434898 548490 435134
rect 548726 434898 548768 435134
rect 548448 434866 548768 434898
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 24114 385774 24734 421218
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 41568 403174 41888 403206
rect 41568 402938 41610 403174
rect 41846 402938 41888 403174
rect 41568 402854 41888 402938
rect 41568 402618 41610 402854
rect 41846 402618 41888 402854
rect 41568 402586 41888 402618
rect 72288 403174 72608 403206
rect 72288 402938 72330 403174
rect 72566 402938 72608 403174
rect 72288 402854 72608 402938
rect 72288 402618 72330 402854
rect 72566 402618 72608 402854
rect 72288 402586 72608 402618
rect 103008 403174 103328 403206
rect 103008 402938 103050 403174
rect 103286 402938 103328 403174
rect 103008 402854 103328 402938
rect 103008 402618 103050 402854
rect 103286 402618 103328 402854
rect 103008 402586 103328 402618
rect 133728 403174 134048 403206
rect 133728 402938 133770 403174
rect 134006 402938 134048 403174
rect 133728 402854 134048 402938
rect 133728 402618 133770 402854
rect 134006 402618 134048 402854
rect 133728 402586 134048 402618
rect 164448 403174 164768 403206
rect 164448 402938 164490 403174
rect 164726 402938 164768 403174
rect 164448 402854 164768 402938
rect 164448 402618 164490 402854
rect 164726 402618 164768 402854
rect 164448 402586 164768 402618
rect 195168 403174 195488 403206
rect 195168 402938 195210 403174
rect 195446 402938 195488 403174
rect 195168 402854 195488 402938
rect 195168 402618 195210 402854
rect 195446 402618 195488 402854
rect 195168 402586 195488 402618
rect 225888 403174 226208 403206
rect 225888 402938 225930 403174
rect 226166 402938 226208 403174
rect 225888 402854 226208 402938
rect 225888 402618 225930 402854
rect 226166 402618 226208 402854
rect 225888 402586 226208 402618
rect 256608 403174 256928 403206
rect 256608 402938 256650 403174
rect 256886 402938 256928 403174
rect 256608 402854 256928 402938
rect 256608 402618 256650 402854
rect 256886 402618 256928 402854
rect 256608 402586 256928 402618
rect 287328 403174 287648 403206
rect 287328 402938 287370 403174
rect 287606 402938 287648 403174
rect 287328 402854 287648 402938
rect 287328 402618 287370 402854
rect 287606 402618 287648 402854
rect 287328 402586 287648 402618
rect 318048 403174 318368 403206
rect 318048 402938 318090 403174
rect 318326 402938 318368 403174
rect 318048 402854 318368 402938
rect 318048 402618 318090 402854
rect 318326 402618 318368 402854
rect 318048 402586 318368 402618
rect 348768 403174 349088 403206
rect 348768 402938 348810 403174
rect 349046 402938 349088 403174
rect 348768 402854 349088 402938
rect 348768 402618 348810 402854
rect 349046 402618 349088 402854
rect 348768 402586 349088 402618
rect 379488 403174 379808 403206
rect 379488 402938 379530 403174
rect 379766 402938 379808 403174
rect 379488 402854 379808 402938
rect 379488 402618 379530 402854
rect 379766 402618 379808 402854
rect 379488 402586 379808 402618
rect 410208 403174 410528 403206
rect 410208 402938 410250 403174
rect 410486 402938 410528 403174
rect 410208 402854 410528 402938
rect 410208 402618 410250 402854
rect 410486 402618 410528 402854
rect 410208 402586 410528 402618
rect 440928 403174 441248 403206
rect 440928 402938 440970 403174
rect 441206 402938 441248 403174
rect 440928 402854 441248 402938
rect 440928 402618 440970 402854
rect 441206 402618 441248 402854
rect 440928 402586 441248 402618
rect 471648 403174 471968 403206
rect 471648 402938 471690 403174
rect 471926 402938 471968 403174
rect 471648 402854 471968 402938
rect 471648 402618 471690 402854
rect 471926 402618 471968 402854
rect 471648 402586 471968 402618
rect 502368 403174 502688 403206
rect 502368 402938 502410 403174
rect 502646 402938 502688 403174
rect 502368 402854 502688 402938
rect 502368 402618 502410 402854
rect 502646 402618 502688 402854
rect 502368 402586 502688 402618
rect 533088 403174 533408 403206
rect 533088 402938 533130 403174
rect 533366 402938 533408 403174
rect 533088 402854 533408 402938
rect 533088 402618 533130 402854
rect 533366 402618 533408 402854
rect 533088 402586 533408 402618
rect 26208 399454 26528 399486
rect 26208 399218 26250 399454
rect 26486 399218 26528 399454
rect 26208 399134 26528 399218
rect 26208 398898 26250 399134
rect 26486 398898 26528 399134
rect 26208 398866 26528 398898
rect 56928 399454 57248 399486
rect 56928 399218 56970 399454
rect 57206 399218 57248 399454
rect 56928 399134 57248 399218
rect 56928 398898 56970 399134
rect 57206 398898 57248 399134
rect 56928 398866 57248 398898
rect 87648 399454 87968 399486
rect 87648 399218 87690 399454
rect 87926 399218 87968 399454
rect 87648 399134 87968 399218
rect 87648 398898 87690 399134
rect 87926 398898 87968 399134
rect 87648 398866 87968 398898
rect 118368 399454 118688 399486
rect 118368 399218 118410 399454
rect 118646 399218 118688 399454
rect 118368 399134 118688 399218
rect 118368 398898 118410 399134
rect 118646 398898 118688 399134
rect 118368 398866 118688 398898
rect 149088 399454 149408 399486
rect 149088 399218 149130 399454
rect 149366 399218 149408 399454
rect 149088 399134 149408 399218
rect 149088 398898 149130 399134
rect 149366 398898 149408 399134
rect 149088 398866 149408 398898
rect 179808 399454 180128 399486
rect 179808 399218 179850 399454
rect 180086 399218 180128 399454
rect 179808 399134 180128 399218
rect 179808 398898 179850 399134
rect 180086 398898 180128 399134
rect 179808 398866 180128 398898
rect 210528 399454 210848 399486
rect 210528 399218 210570 399454
rect 210806 399218 210848 399454
rect 210528 399134 210848 399218
rect 210528 398898 210570 399134
rect 210806 398898 210848 399134
rect 210528 398866 210848 398898
rect 241248 399454 241568 399486
rect 241248 399218 241290 399454
rect 241526 399218 241568 399454
rect 241248 399134 241568 399218
rect 241248 398898 241290 399134
rect 241526 398898 241568 399134
rect 241248 398866 241568 398898
rect 271968 399454 272288 399486
rect 271968 399218 272010 399454
rect 272246 399218 272288 399454
rect 271968 399134 272288 399218
rect 271968 398898 272010 399134
rect 272246 398898 272288 399134
rect 271968 398866 272288 398898
rect 302688 399454 303008 399486
rect 302688 399218 302730 399454
rect 302966 399218 303008 399454
rect 302688 399134 303008 399218
rect 302688 398898 302730 399134
rect 302966 398898 303008 399134
rect 302688 398866 303008 398898
rect 333408 399454 333728 399486
rect 333408 399218 333450 399454
rect 333686 399218 333728 399454
rect 333408 399134 333728 399218
rect 333408 398898 333450 399134
rect 333686 398898 333728 399134
rect 333408 398866 333728 398898
rect 364128 399454 364448 399486
rect 364128 399218 364170 399454
rect 364406 399218 364448 399454
rect 364128 399134 364448 399218
rect 364128 398898 364170 399134
rect 364406 398898 364448 399134
rect 364128 398866 364448 398898
rect 394848 399454 395168 399486
rect 394848 399218 394890 399454
rect 395126 399218 395168 399454
rect 394848 399134 395168 399218
rect 394848 398898 394890 399134
rect 395126 398898 395168 399134
rect 394848 398866 395168 398898
rect 425568 399454 425888 399486
rect 425568 399218 425610 399454
rect 425846 399218 425888 399454
rect 425568 399134 425888 399218
rect 425568 398898 425610 399134
rect 425846 398898 425888 399134
rect 425568 398866 425888 398898
rect 456288 399454 456608 399486
rect 456288 399218 456330 399454
rect 456566 399218 456608 399454
rect 456288 399134 456608 399218
rect 456288 398898 456330 399134
rect 456566 398898 456608 399134
rect 456288 398866 456608 398898
rect 487008 399454 487328 399486
rect 487008 399218 487050 399454
rect 487286 399218 487328 399454
rect 487008 399134 487328 399218
rect 487008 398898 487050 399134
rect 487286 398898 487328 399134
rect 487008 398866 487328 398898
rect 517728 399454 518048 399486
rect 517728 399218 517770 399454
rect 518006 399218 518048 399454
rect 517728 399134 518048 399218
rect 517728 398898 517770 399134
rect 518006 398898 518048 399134
rect 517728 398866 518048 398898
rect 548448 399454 548768 399486
rect 548448 399218 548490 399454
rect 548726 399218 548768 399454
rect 548448 399134 548768 399218
rect 548448 398898 548490 399134
rect 548726 398898 548768 399134
rect 548448 398866 548768 398898
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 24114 349774 24734 385218
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 41568 367174 41888 367206
rect 41568 366938 41610 367174
rect 41846 366938 41888 367174
rect 41568 366854 41888 366938
rect 41568 366618 41610 366854
rect 41846 366618 41888 366854
rect 41568 366586 41888 366618
rect 72288 367174 72608 367206
rect 72288 366938 72330 367174
rect 72566 366938 72608 367174
rect 72288 366854 72608 366938
rect 72288 366618 72330 366854
rect 72566 366618 72608 366854
rect 72288 366586 72608 366618
rect 103008 367174 103328 367206
rect 103008 366938 103050 367174
rect 103286 366938 103328 367174
rect 103008 366854 103328 366938
rect 103008 366618 103050 366854
rect 103286 366618 103328 366854
rect 103008 366586 103328 366618
rect 133728 367174 134048 367206
rect 133728 366938 133770 367174
rect 134006 366938 134048 367174
rect 133728 366854 134048 366938
rect 133728 366618 133770 366854
rect 134006 366618 134048 366854
rect 133728 366586 134048 366618
rect 164448 367174 164768 367206
rect 164448 366938 164490 367174
rect 164726 366938 164768 367174
rect 164448 366854 164768 366938
rect 164448 366618 164490 366854
rect 164726 366618 164768 366854
rect 164448 366586 164768 366618
rect 195168 367174 195488 367206
rect 195168 366938 195210 367174
rect 195446 366938 195488 367174
rect 195168 366854 195488 366938
rect 195168 366618 195210 366854
rect 195446 366618 195488 366854
rect 195168 366586 195488 366618
rect 225888 367174 226208 367206
rect 225888 366938 225930 367174
rect 226166 366938 226208 367174
rect 225888 366854 226208 366938
rect 225888 366618 225930 366854
rect 226166 366618 226208 366854
rect 225888 366586 226208 366618
rect 256608 367174 256928 367206
rect 256608 366938 256650 367174
rect 256886 366938 256928 367174
rect 256608 366854 256928 366938
rect 256608 366618 256650 366854
rect 256886 366618 256928 366854
rect 256608 366586 256928 366618
rect 287328 367174 287648 367206
rect 287328 366938 287370 367174
rect 287606 366938 287648 367174
rect 287328 366854 287648 366938
rect 287328 366618 287370 366854
rect 287606 366618 287648 366854
rect 287328 366586 287648 366618
rect 318048 367174 318368 367206
rect 318048 366938 318090 367174
rect 318326 366938 318368 367174
rect 318048 366854 318368 366938
rect 318048 366618 318090 366854
rect 318326 366618 318368 366854
rect 318048 366586 318368 366618
rect 348768 367174 349088 367206
rect 348768 366938 348810 367174
rect 349046 366938 349088 367174
rect 348768 366854 349088 366938
rect 348768 366618 348810 366854
rect 349046 366618 349088 366854
rect 348768 366586 349088 366618
rect 379488 367174 379808 367206
rect 379488 366938 379530 367174
rect 379766 366938 379808 367174
rect 379488 366854 379808 366938
rect 379488 366618 379530 366854
rect 379766 366618 379808 366854
rect 379488 366586 379808 366618
rect 410208 367174 410528 367206
rect 410208 366938 410250 367174
rect 410486 366938 410528 367174
rect 410208 366854 410528 366938
rect 410208 366618 410250 366854
rect 410486 366618 410528 366854
rect 410208 366586 410528 366618
rect 440928 367174 441248 367206
rect 440928 366938 440970 367174
rect 441206 366938 441248 367174
rect 440928 366854 441248 366938
rect 440928 366618 440970 366854
rect 441206 366618 441248 366854
rect 440928 366586 441248 366618
rect 471648 367174 471968 367206
rect 471648 366938 471690 367174
rect 471926 366938 471968 367174
rect 471648 366854 471968 366938
rect 471648 366618 471690 366854
rect 471926 366618 471968 366854
rect 471648 366586 471968 366618
rect 502368 367174 502688 367206
rect 502368 366938 502410 367174
rect 502646 366938 502688 367174
rect 502368 366854 502688 366938
rect 502368 366618 502410 366854
rect 502646 366618 502688 366854
rect 502368 366586 502688 366618
rect 533088 367174 533408 367206
rect 533088 366938 533130 367174
rect 533366 366938 533408 367174
rect 533088 366854 533408 366938
rect 533088 366618 533130 366854
rect 533366 366618 533408 366854
rect 533088 366586 533408 366618
rect 26208 363454 26528 363486
rect 26208 363218 26250 363454
rect 26486 363218 26528 363454
rect 26208 363134 26528 363218
rect 26208 362898 26250 363134
rect 26486 362898 26528 363134
rect 26208 362866 26528 362898
rect 56928 363454 57248 363486
rect 56928 363218 56970 363454
rect 57206 363218 57248 363454
rect 56928 363134 57248 363218
rect 56928 362898 56970 363134
rect 57206 362898 57248 363134
rect 56928 362866 57248 362898
rect 87648 363454 87968 363486
rect 87648 363218 87690 363454
rect 87926 363218 87968 363454
rect 87648 363134 87968 363218
rect 87648 362898 87690 363134
rect 87926 362898 87968 363134
rect 87648 362866 87968 362898
rect 118368 363454 118688 363486
rect 118368 363218 118410 363454
rect 118646 363218 118688 363454
rect 118368 363134 118688 363218
rect 118368 362898 118410 363134
rect 118646 362898 118688 363134
rect 118368 362866 118688 362898
rect 149088 363454 149408 363486
rect 149088 363218 149130 363454
rect 149366 363218 149408 363454
rect 149088 363134 149408 363218
rect 149088 362898 149130 363134
rect 149366 362898 149408 363134
rect 149088 362866 149408 362898
rect 179808 363454 180128 363486
rect 179808 363218 179850 363454
rect 180086 363218 180128 363454
rect 179808 363134 180128 363218
rect 179808 362898 179850 363134
rect 180086 362898 180128 363134
rect 179808 362866 180128 362898
rect 210528 363454 210848 363486
rect 210528 363218 210570 363454
rect 210806 363218 210848 363454
rect 210528 363134 210848 363218
rect 210528 362898 210570 363134
rect 210806 362898 210848 363134
rect 210528 362866 210848 362898
rect 241248 363454 241568 363486
rect 241248 363218 241290 363454
rect 241526 363218 241568 363454
rect 241248 363134 241568 363218
rect 241248 362898 241290 363134
rect 241526 362898 241568 363134
rect 241248 362866 241568 362898
rect 271968 363454 272288 363486
rect 271968 363218 272010 363454
rect 272246 363218 272288 363454
rect 271968 363134 272288 363218
rect 271968 362898 272010 363134
rect 272246 362898 272288 363134
rect 271968 362866 272288 362898
rect 302688 363454 303008 363486
rect 302688 363218 302730 363454
rect 302966 363218 303008 363454
rect 302688 363134 303008 363218
rect 302688 362898 302730 363134
rect 302966 362898 303008 363134
rect 302688 362866 303008 362898
rect 333408 363454 333728 363486
rect 333408 363218 333450 363454
rect 333686 363218 333728 363454
rect 333408 363134 333728 363218
rect 333408 362898 333450 363134
rect 333686 362898 333728 363134
rect 333408 362866 333728 362898
rect 364128 363454 364448 363486
rect 364128 363218 364170 363454
rect 364406 363218 364448 363454
rect 364128 363134 364448 363218
rect 364128 362898 364170 363134
rect 364406 362898 364448 363134
rect 364128 362866 364448 362898
rect 394848 363454 395168 363486
rect 394848 363218 394890 363454
rect 395126 363218 395168 363454
rect 394848 363134 395168 363218
rect 394848 362898 394890 363134
rect 395126 362898 395168 363134
rect 394848 362866 395168 362898
rect 425568 363454 425888 363486
rect 425568 363218 425610 363454
rect 425846 363218 425888 363454
rect 425568 363134 425888 363218
rect 425568 362898 425610 363134
rect 425846 362898 425888 363134
rect 425568 362866 425888 362898
rect 456288 363454 456608 363486
rect 456288 363218 456330 363454
rect 456566 363218 456608 363454
rect 456288 363134 456608 363218
rect 456288 362898 456330 363134
rect 456566 362898 456608 363134
rect 456288 362866 456608 362898
rect 487008 363454 487328 363486
rect 487008 363218 487050 363454
rect 487286 363218 487328 363454
rect 487008 363134 487328 363218
rect 487008 362898 487050 363134
rect 487286 362898 487328 363134
rect 487008 362866 487328 362898
rect 517728 363454 518048 363486
rect 517728 363218 517770 363454
rect 518006 363218 518048 363454
rect 517728 363134 518048 363218
rect 517728 362898 517770 363134
rect 518006 362898 518048 363134
rect 517728 362866 518048 362898
rect 548448 363454 548768 363486
rect 548448 363218 548490 363454
rect 548726 363218 548768 363454
rect 548448 363134 548768 363218
rect 548448 362898 548490 363134
rect 548726 362898 548768 363134
rect 548448 362866 548768 362898
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 24114 313774 24734 349218
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 41568 331174 41888 331206
rect 41568 330938 41610 331174
rect 41846 330938 41888 331174
rect 41568 330854 41888 330938
rect 41568 330618 41610 330854
rect 41846 330618 41888 330854
rect 41568 330586 41888 330618
rect 72288 331174 72608 331206
rect 72288 330938 72330 331174
rect 72566 330938 72608 331174
rect 72288 330854 72608 330938
rect 72288 330618 72330 330854
rect 72566 330618 72608 330854
rect 72288 330586 72608 330618
rect 103008 331174 103328 331206
rect 103008 330938 103050 331174
rect 103286 330938 103328 331174
rect 103008 330854 103328 330938
rect 103008 330618 103050 330854
rect 103286 330618 103328 330854
rect 103008 330586 103328 330618
rect 133728 331174 134048 331206
rect 133728 330938 133770 331174
rect 134006 330938 134048 331174
rect 133728 330854 134048 330938
rect 133728 330618 133770 330854
rect 134006 330618 134048 330854
rect 133728 330586 134048 330618
rect 164448 331174 164768 331206
rect 164448 330938 164490 331174
rect 164726 330938 164768 331174
rect 164448 330854 164768 330938
rect 164448 330618 164490 330854
rect 164726 330618 164768 330854
rect 164448 330586 164768 330618
rect 195168 331174 195488 331206
rect 195168 330938 195210 331174
rect 195446 330938 195488 331174
rect 195168 330854 195488 330938
rect 195168 330618 195210 330854
rect 195446 330618 195488 330854
rect 195168 330586 195488 330618
rect 225888 331174 226208 331206
rect 225888 330938 225930 331174
rect 226166 330938 226208 331174
rect 225888 330854 226208 330938
rect 225888 330618 225930 330854
rect 226166 330618 226208 330854
rect 225888 330586 226208 330618
rect 256608 331174 256928 331206
rect 256608 330938 256650 331174
rect 256886 330938 256928 331174
rect 256608 330854 256928 330938
rect 256608 330618 256650 330854
rect 256886 330618 256928 330854
rect 256608 330586 256928 330618
rect 287328 331174 287648 331206
rect 287328 330938 287370 331174
rect 287606 330938 287648 331174
rect 287328 330854 287648 330938
rect 287328 330618 287370 330854
rect 287606 330618 287648 330854
rect 287328 330586 287648 330618
rect 318048 331174 318368 331206
rect 318048 330938 318090 331174
rect 318326 330938 318368 331174
rect 318048 330854 318368 330938
rect 318048 330618 318090 330854
rect 318326 330618 318368 330854
rect 318048 330586 318368 330618
rect 348768 331174 349088 331206
rect 348768 330938 348810 331174
rect 349046 330938 349088 331174
rect 348768 330854 349088 330938
rect 348768 330618 348810 330854
rect 349046 330618 349088 330854
rect 348768 330586 349088 330618
rect 379488 331174 379808 331206
rect 379488 330938 379530 331174
rect 379766 330938 379808 331174
rect 379488 330854 379808 330938
rect 379488 330618 379530 330854
rect 379766 330618 379808 330854
rect 379488 330586 379808 330618
rect 410208 331174 410528 331206
rect 410208 330938 410250 331174
rect 410486 330938 410528 331174
rect 410208 330854 410528 330938
rect 410208 330618 410250 330854
rect 410486 330618 410528 330854
rect 410208 330586 410528 330618
rect 440928 331174 441248 331206
rect 440928 330938 440970 331174
rect 441206 330938 441248 331174
rect 440928 330854 441248 330938
rect 440928 330618 440970 330854
rect 441206 330618 441248 330854
rect 440928 330586 441248 330618
rect 471648 331174 471968 331206
rect 471648 330938 471690 331174
rect 471926 330938 471968 331174
rect 471648 330854 471968 330938
rect 471648 330618 471690 330854
rect 471926 330618 471968 330854
rect 471648 330586 471968 330618
rect 502368 331174 502688 331206
rect 502368 330938 502410 331174
rect 502646 330938 502688 331174
rect 502368 330854 502688 330938
rect 502368 330618 502410 330854
rect 502646 330618 502688 330854
rect 502368 330586 502688 330618
rect 533088 331174 533408 331206
rect 533088 330938 533130 331174
rect 533366 330938 533408 331174
rect 533088 330854 533408 330938
rect 533088 330618 533130 330854
rect 533366 330618 533408 330854
rect 533088 330586 533408 330618
rect 26208 327454 26528 327486
rect 26208 327218 26250 327454
rect 26486 327218 26528 327454
rect 26208 327134 26528 327218
rect 26208 326898 26250 327134
rect 26486 326898 26528 327134
rect 26208 326866 26528 326898
rect 56928 327454 57248 327486
rect 56928 327218 56970 327454
rect 57206 327218 57248 327454
rect 56928 327134 57248 327218
rect 56928 326898 56970 327134
rect 57206 326898 57248 327134
rect 56928 326866 57248 326898
rect 87648 327454 87968 327486
rect 87648 327218 87690 327454
rect 87926 327218 87968 327454
rect 87648 327134 87968 327218
rect 87648 326898 87690 327134
rect 87926 326898 87968 327134
rect 87648 326866 87968 326898
rect 118368 327454 118688 327486
rect 118368 327218 118410 327454
rect 118646 327218 118688 327454
rect 118368 327134 118688 327218
rect 118368 326898 118410 327134
rect 118646 326898 118688 327134
rect 118368 326866 118688 326898
rect 149088 327454 149408 327486
rect 149088 327218 149130 327454
rect 149366 327218 149408 327454
rect 149088 327134 149408 327218
rect 149088 326898 149130 327134
rect 149366 326898 149408 327134
rect 149088 326866 149408 326898
rect 179808 327454 180128 327486
rect 179808 327218 179850 327454
rect 180086 327218 180128 327454
rect 179808 327134 180128 327218
rect 179808 326898 179850 327134
rect 180086 326898 180128 327134
rect 179808 326866 180128 326898
rect 210528 327454 210848 327486
rect 210528 327218 210570 327454
rect 210806 327218 210848 327454
rect 210528 327134 210848 327218
rect 210528 326898 210570 327134
rect 210806 326898 210848 327134
rect 210528 326866 210848 326898
rect 241248 327454 241568 327486
rect 241248 327218 241290 327454
rect 241526 327218 241568 327454
rect 241248 327134 241568 327218
rect 241248 326898 241290 327134
rect 241526 326898 241568 327134
rect 241248 326866 241568 326898
rect 271968 327454 272288 327486
rect 271968 327218 272010 327454
rect 272246 327218 272288 327454
rect 271968 327134 272288 327218
rect 271968 326898 272010 327134
rect 272246 326898 272288 327134
rect 271968 326866 272288 326898
rect 302688 327454 303008 327486
rect 302688 327218 302730 327454
rect 302966 327218 303008 327454
rect 302688 327134 303008 327218
rect 302688 326898 302730 327134
rect 302966 326898 303008 327134
rect 302688 326866 303008 326898
rect 333408 327454 333728 327486
rect 333408 327218 333450 327454
rect 333686 327218 333728 327454
rect 333408 327134 333728 327218
rect 333408 326898 333450 327134
rect 333686 326898 333728 327134
rect 333408 326866 333728 326898
rect 364128 327454 364448 327486
rect 364128 327218 364170 327454
rect 364406 327218 364448 327454
rect 364128 327134 364448 327218
rect 364128 326898 364170 327134
rect 364406 326898 364448 327134
rect 364128 326866 364448 326898
rect 394848 327454 395168 327486
rect 394848 327218 394890 327454
rect 395126 327218 395168 327454
rect 394848 327134 395168 327218
rect 394848 326898 394890 327134
rect 395126 326898 395168 327134
rect 394848 326866 395168 326898
rect 425568 327454 425888 327486
rect 425568 327218 425610 327454
rect 425846 327218 425888 327454
rect 425568 327134 425888 327218
rect 425568 326898 425610 327134
rect 425846 326898 425888 327134
rect 425568 326866 425888 326898
rect 456288 327454 456608 327486
rect 456288 327218 456330 327454
rect 456566 327218 456608 327454
rect 456288 327134 456608 327218
rect 456288 326898 456330 327134
rect 456566 326898 456608 327134
rect 456288 326866 456608 326898
rect 487008 327454 487328 327486
rect 487008 327218 487050 327454
rect 487286 327218 487328 327454
rect 487008 327134 487328 327218
rect 487008 326898 487050 327134
rect 487286 326898 487328 327134
rect 487008 326866 487328 326898
rect 517728 327454 518048 327486
rect 517728 327218 517770 327454
rect 518006 327218 518048 327454
rect 517728 327134 518048 327218
rect 517728 326898 517770 327134
rect 518006 326898 518048 327134
rect 517728 326866 518048 326898
rect 548448 327454 548768 327486
rect 548448 327218 548490 327454
rect 548726 327218 548768 327454
rect 548448 327134 548768 327218
rect 548448 326898 548490 327134
rect 548726 326898 548768 327134
rect 548448 326866 548768 326898
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 24114 277774 24734 313218
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 41568 295174 41888 295206
rect 41568 294938 41610 295174
rect 41846 294938 41888 295174
rect 41568 294854 41888 294938
rect 41568 294618 41610 294854
rect 41846 294618 41888 294854
rect 41568 294586 41888 294618
rect 72288 295174 72608 295206
rect 72288 294938 72330 295174
rect 72566 294938 72608 295174
rect 72288 294854 72608 294938
rect 72288 294618 72330 294854
rect 72566 294618 72608 294854
rect 72288 294586 72608 294618
rect 103008 295174 103328 295206
rect 103008 294938 103050 295174
rect 103286 294938 103328 295174
rect 103008 294854 103328 294938
rect 103008 294618 103050 294854
rect 103286 294618 103328 294854
rect 103008 294586 103328 294618
rect 133728 295174 134048 295206
rect 133728 294938 133770 295174
rect 134006 294938 134048 295174
rect 133728 294854 134048 294938
rect 133728 294618 133770 294854
rect 134006 294618 134048 294854
rect 133728 294586 134048 294618
rect 164448 295174 164768 295206
rect 164448 294938 164490 295174
rect 164726 294938 164768 295174
rect 164448 294854 164768 294938
rect 164448 294618 164490 294854
rect 164726 294618 164768 294854
rect 164448 294586 164768 294618
rect 195168 295174 195488 295206
rect 195168 294938 195210 295174
rect 195446 294938 195488 295174
rect 195168 294854 195488 294938
rect 195168 294618 195210 294854
rect 195446 294618 195488 294854
rect 195168 294586 195488 294618
rect 225888 295174 226208 295206
rect 225888 294938 225930 295174
rect 226166 294938 226208 295174
rect 225888 294854 226208 294938
rect 225888 294618 225930 294854
rect 226166 294618 226208 294854
rect 225888 294586 226208 294618
rect 256608 295174 256928 295206
rect 256608 294938 256650 295174
rect 256886 294938 256928 295174
rect 256608 294854 256928 294938
rect 256608 294618 256650 294854
rect 256886 294618 256928 294854
rect 256608 294586 256928 294618
rect 287328 295174 287648 295206
rect 287328 294938 287370 295174
rect 287606 294938 287648 295174
rect 287328 294854 287648 294938
rect 287328 294618 287370 294854
rect 287606 294618 287648 294854
rect 287328 294586 287648 294618
rect 318048 295174 318368 295206
rect 318048 294938 318090 295174
rect 318326 294938 318368 295174
rect 318048 294854 318368 294938
rect 318048 294618 318090 294854
rect 318326 294618 318368 294854
rect 318048 294586 318368 294618
rect 348768 295174 349088 295206
rect 348768 294938 348810 295174
rect 349046 294938 349088 295174
rect 348768 294854 349088 294938
rect 348768 294618 348810 294854
rect 349046 294618 349088 294854
rect 348768 294586 349088 294618
rect 379488 295174 379808 295206
rect 379488 294938 379530 295174
rect 379766 294938 379808 295174
rect 379488 294854 379808 294938
rect 379488 294618 379530 294854
rect 379766 294618 379808 294854
rect 379488 294586 379808 294618
rect 410208 295174 410528 295206
rect 410208 294938 410250 295174
rect 410486 294938 410528 295174
rect 410208 294854 410528 294938
rect 410208 294618 410250 294854
rect 410486 294618 410528 294854
rect 410208 294586 410528 294618
rect 440928 295174 441248 295206
rect 440928 294938 440970 295174
rect 441206 294938 441248 295174
rect 440928 294854 441248 294938
rect 440928 294618 440970 294854
rect 441206 294618 441248 294854
rect 440928 294586 441248 294618
rect 471648 295174 471968 295206
rect 471648 294938 471690 295174
rect 471926 294938 471968 295174
rect 471648 294854 471968 294938
rect 471648 294618 471690 294854
rect 471926 294618 471968 294854
rect 471648 294586 471968 294618
rect 502368 295174 502688 295206
rect 502368 294938 502410 295174
rect 502646 294938 502688 295174
rect 502368 294854 502688 294938
rect 502368 294618 502410 294854
rect 502646 294618 502688 294854
rect 502368 294586 502688 294618
rect 533088 295174 533408 295206
rect 533088 294938 533130 295174
rect 533366 294938 533408 295174
rect 533088 294854 533408 294938
rect 533088 294618 533130 294854
rect 533366 294618 533408 294854
rect 533088 294586 533408 294618
rect 26208 291454 26528 291486
rect 26208 291218 26250 291454
rect 26486 291218 26528 291454
rect 26208 291134 26528 291218
rect 26208 290898 26250 291134
rect 26486 290898 26528 291134
rect 26208 290866 26528 290898
rect 56928 291454 57248 291486
rect 56928 291218 56970 291454
rect 57206 291218 57248 291454
rect 56928 291134 57248 291218
rect 56928 290898 56970 291134
rect 57206 290898 57248 291134
rect 56928 290866 57248 290898
rect 87648 291454 87968 291486
rect 87648 291218 87690 291454
rect 87926 291218 87968 291454
rect 87648 291134 87968 291218
rect 87648 290898 87690 291134
rect 87926 290898 87968 291134
rect 87648 290866 87968 290898
rect 118368 291454 118688 291486
rect 118368 291218 118410 291454
rect 118646 291218 118688 291454
rect 118368 291134 118688 291218
rect 118368 290898 118410 291134
rect 118646 290898 118688 291134
rect 118368 290866 118688 290898
rect 149088 291454 149408 291486
rect 149088 291218 149130 291454
rect 149366 291218 149408 291454
rect 149088 291134 149408 291218
rect 149088 290898 149130 291134
rect 149366 290898 149408 291134
rect 149088 290866 149408 290898
rect 179808 291454 180128 291486
rect 179808 291218 179850 291454
rect 180086 291218 180128 291454
rect 179808 291134 180128 291218
rect 179808 290898 179850 291134
rect 180086 290898 180128 291134
rect 179808 290866 180128 290898
rect 210528 291454 210848 291486
rect 210528 291218 210570 291454
rect 210806 291218 210848 291454
rect 210528 291134 210848 291218
rect 210528 290898 210570 291134
rect 210806 290898 210848 291134
rect 210528 290866 210848 290898
rect 241248 291454 241568 291486
rect 241248 291218 241290 291454
rect 241526 291218 241568 291454
rect 241248 291134 241568 291218
rect 241248 290898 241290 291134
rect 241526 290898 241568 291134
rect 241248 290866 241568 290898
rect 271968 291454 272288 291486
rect 271968 291218 272010 291454
rect 272246 291218 272288 291454
rect 271968 291134 272288 291218
rect 271968 290898 272010 291134
rect 272246 290898 272288 291134
rect 271968 290866 272288 290898
rect 302688 291454 303008 291486
rect 302688 291218 302730 291454
rect 302966 291218 303008 291454
rect 302688 291134 303008 291218
rect 302688 290898 302730 291134
rect 302966 290898 303008 291134
rect 302688 290866 303008 290898
rect 333408 291454 333728 291486
rect 333408 291218 333450 291454
rect 333686 291218 333728 291454
rect 333408 291134 333728 291218
rect 333408 290898 333450 291134
rect 333686 290898 333728 291134
rect 333408 290866 333728 290898
rect 364128 291454 364448 291486
rect 364128 291218 364170 291454
rect 364406 291218 364448 291454
rect 364128 291134 364448 291218
rect 364128 290898 364170 291134
rect 364406 290898 364448 291134
rect 364128 290866 364448 290898
rect 394848 291454 395168 291486
rect 394848 291218 394890 291454
rect 395126 291218 395168 291454
rect 394848 291134 395168 291218
rect 394848 290898 394890 291134
rect 395126 290898 395168 291134
rect 394848 290866 395168 290898
rect 425568 291454 425888 291486
rect 425568 291218 425610 291454
rect 425846 291218 425888 291454
rect 425568 291134 425888 291218
rect 425568 290898 425610 291134
rect 425846 290898 425888 291134
rect 425568 290866 425888 290898
rect 456288 291454 456608 291486
rect 456288 291218 456330 291454
rect 456566 291218 456608 291454
rect 456288 291134 456608 291218
rect 456288 290898 456330 291134
rect 456566 290898 456608 291134
rect 456288 290866 456608 290898
rect 487008 291454 487328 291486
rect 487008 291218 487050 291454
rect 487286 291218 487328 291454
rect 487008 291134 487328 291218
rect 487008 290898 487050 291134
rect 487286 290898 487328 291134
rect 487008 290866 487328 290898
rect 517728 291454 518048 291486
rect 517728 291218 517770 291454
rect 518006 291218 518048 291454
rect 517728 291134 518048 291218
rect 517728 290898 517770 291134
rect 518006 290898 518048 291134
rect 517728 290866 518048 290898
rect 548448 291454 548768 291486
rect 548448 291218 548490 291454
rect 548726 291218 548768 291454
rect 548448 291134 548768 291218
rect 548448 290898 548490 291134
rect 548726 290898 548768 291134
rect 548448 290866 548768 290898
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 24114 241774 24734 277218
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 41568 259174 41888 259206
rect 41568 258938 41610 259174
rect 41846 258938 41888 259174
rect 41568 258854 41888 258938
rect 41568 258618 41610 258854
rect 41846 258618 41888 258854
rect 41568 258586 41888 258618
rect 72288 259174 72608 259206
rect 72288 258938 72330 259174
rect 72566 258938 72608 259174
rect 72288 258854 72608 258938
rect 72288 258618 72330 258854
rect 72566 258618 72608 258854
rect 72288 258586 72608 258618
rect 103008 259174 103328 259206
rect 103008 258938 103050 259174
rect 103286 258938 103328 259174
rect 103008 258854 103328 258938
rect 103008 258618 103050 258854
rect 103286 258618 103328 258854
rect 103008 258586 103328 258618
rect 133728 259174 134048 259206
rect 133728 258938 133770 259174
rect 134006 258938 134048 259174
rect 133728 258854 134048 258938
rect 133728 258618 133770 258854
rect 134006 258618 134048 258854
rect 133728 258586 134048 258618
rect 164448 259174 164768 259206
rect 164448 258938 164490 259174
rect 164726 258938 164768 259174
rect 164448 258854 164768 258938
rect 164448 258618 164490 258854
rect 164726 258618 164768 258854
rect 164448 258586 164768 258618
rect 195168 259174 195488 259206
rect 195168 258938 195210 259174
rect 195446 258938 195488 259174
rect 195168 258854 195488 258938
rect 195168 258618 195210 258854
rect 195446 258618 195488 258854
rect 195168 258586 195488 258618
rect 225888 259174 226208 259206
rect 225888 258938 225930 259174
rect 226166 258938 226208 259174
rect 225888 258854 226208 258938
rect 225888 258618 225930 258854
rect 226166 258618 226208 258854
rect 225888 258586 226208 258618
rect 256608 259174 256928 259206
rect 256608 258938 256650 259174
rect 256886 258938 256928 259174
rect 256608 258854 256928 258938
rect 256608 258618 256650 258854
rect 256886 258618 256928 258854
rect 256608 258586 256928 258618
rect 287328 259174 287648 259206
rect 287328 258938 287370 259174
rect 287606 258938 287648 259174
rect 287328 258854 287648 258938
rect 287328 258618 287370 258854
rect 287606 258618 287648 258854
rect 287328 258586 287648 258618
rect 318048 259174 318368 259206
rect 318048 258938 318090 259174
rect 318326 258938 318368 259174
rect 318048 258854 318368 258938
rect 318048 258618 318090 258854
rect 318326 258618 318368 258854
rect 318048 258586 318368 258618
rect 348768 259174 349088 259206
rect 348768 258938 348810 259174
rect 349046 258938 349088 259174
rect 348768 258854 349088 258938
rect 348768 258618 348810 258854
rect 349046 258618 349088 258854
rect 348768 258586 349088 258618
rect 379488 259174 379808 259206
rect 379488 258938 379530 259174
rect 379766 258938 379808 259174
rect 379488 258854 379808 258938
rect 379488 258618 379530 258854
rect 379766 258618 379808 258854
rect 379488 258586 379808 258618
rect 410208 259174 410528 259206
rect 410208 258938 410250 259174
rect 410486 258938 410528 259174
rect 410208 258854 410528 258938
rect 410208 258618 410250 258854
rect 410486 258618 410528 258854
rect 410208 258586 410528 258618
rect 440928 259174 441248 259206
rect 440928 258938 440970 259174
rect 441206 258938 441248 259174
rect 440928 258854 441248 258938
rect 440928 258618 440970 258854
rect 441206 258618 441248 258854
rect 440928 258586 441248 258618
rect 471648 259174 471968 259206
rect 471648 258938 471690 259174
rect 471926 258938 471968 259174
rect 471648 258854 471968 258938
rect 471648 258618 471690 258854
rect 471926 258618 471968 258854
rect 471648 258586 471968 258618
rect 502368 259174 502688 259206
rect 502368 258938 502410 259174
rect 502646 258938 502688 259174
rect 502368 258854 502688 258938
rect 502368 258618 502410 258854
rect 502646 258618 502688 258854
rect 502368 258586 502688 258618
rect 533088 259174 533408 259206
rect 533088 258938 533130 259174
rect 533366 258938 533408 259174
rect 533088 258854 533408 258938
rect 533088 258618 533130 258854
rect 533366 258618 533408 258854
rect 533088 258586 533408 258618
rect 26208 255454 26528 255486
rect 26208 255218 26250 255454
rect 26486 255218 26528 255454
rect 26208 255134 26528 255218
rect 26208 254898 26250 255134
rect 26486 254898 26528 255134
rect 26208 254866 26528 254898
rect 56928 255454 57248 255486
rect 56928 255218 56970 255454
rect 57206 255218 57248 255454
rect 56928 255134 57248 255218
rect 56928 254898 56970 255134
rect 57206 254898 57248 255134
rect 56928 254866 57248 254898
rect 87648 255454 87968 255486
rect 87648 255218 87690 255454
rect 87926 255218 87968 255454
rect 87648 255134 87968 255218
rect 87648 254898 87690 255134
rect 87926 254898 87968 255134
rect 87648 254866 87968 254898
rect 118368 255454 118688 255486
rect 118368 255218 118410 255454
rect 118646 255218 118688 255454
rect 118368 255134 118688 255218
rect 118368 254898 118410 255134
rect 118646 254898 118688 255134
rect 118368 254866 118688 254898
rect 149088 255454 149408 255486
rect 149088 255218 149130 255454
rect 149366 255218 149408 255454
rect 149088 255134 149408 255218
rect 149088 254898 149130 255134
rect 149366 254898 149408 255134
rect 149088 254866 149408 254898
rect 179808 255454 180128 255486
rect 179808 255218 179850 255454
rect 180086 255218 180128 255454
rect 179808 255134 180128 255218
rect 179808 254898 179850 255134
rect 180086 254898 180128 255134
rect 179808 254866 180128 254898
rect 210528 255454 210848 255486
rect 210528 255218 210570 255454
rect 210806 255218 210848 255454
rect 210528 255134 210848 255218
rect 210528 254898 210570 255134
rect 210806 254898 210848 255134
rect 210528 254866 210848 254898
rect 241248 255454 241568 255486
rect 241248 255218 241290 255454
rect 241526 255218 241568 255454
rect 241248 255134 241568 255218
rect 241248 254898 241290 255134
rect 241526 254898 241568 255134
rect 241248 254866 241568 254898
rect 271968 255454 272288 255486
rect 271968 255218 272010 255454
rect 272246 255218 272288 255454
rect 271968 255134 272288 255218
rect 271968 254898 272010 255134
rect 272246 254898 272288 255134
rect 271968 254866 272288 254898
rect 302688 255454 303008 255486
rect 302688 255218 302730 255454
rect 302966 255218 303008 255454
rect 302688 255134 303008 255218
rect 302688 254898 302730 255134
rect 302966 254898 303008 255134
rect 302688 254866 303008 254898
rect 333408 255454 333728 255486
rect 333408 255218 333450 255454
rect 333686 255218 333728 255454
rect 333408 255134 333728 255218
rect 333408 254898 333450 255134
rect 333686 254898 333728 255134
rect 333408 254866 333728 254898
rect 364128 255454 364448 255486
rect 364128 255218 364170 255454
rect 364406 255218 364448 255454
rect 364128 255134 364448 255218
rect 364128 254898 364170 255134
rect 364406 254898 364448 255134
rect 364128 254866 364448 254898
rect 394848 255454 395168 255486
rect 394848 255218 394890 255454
rect 395126 255218 395168 255454
rect 394848 255134 395168 255218
rect 394848 254898 394890 255134
rect 395126 254898 395168 255134
rect 394848 254866 395168 254898
rect 425568 255454 425888 255486
rect 425568 255218 425610 255454
rect 425846 255218 425888 255454
rect 425568 255134 425888 255218
rect 425568 254898 425610 255134
rect 425846 254898 425888 255134
rect 425568 254866 425888 254898
rect 456288 255454 456608 255486
rect 456288 255218 456330 255454
rect 456566 255218 456608 255454
rect 456288 255134 456608 255218
rect 456288 254898 456330 255134
rect 456566 254898 456608 255134
rect 456288 254866 456608 254898
rect 487008 255454 487328 255486
rect 487008 255218 487050 255454
rect 487286 255218 487328 255454
rect 487008 255134 487328 255218
rect 487008 254898 487050 255134
rect 487286 254898 487328 255134
rect 487008 254866 487328 254898
rect 517728 255454 518048 255486
rect 517728 255218 517770 255454
rect 518006 255218 518048 255454
rect 517728 255134 518048 255218
rect 517728 254898 517770 255134
rect 518006 254898 518048 255134
rect 517728 254866 518048 254898
rect 548448 255454 548768 255486
rect 548448 255218 548490 255454
rect 548726 255218 548768 255454
rect 548448 255134 548768 255218
rect 548448 254898 548490 255134
rect 548726 254898 548768 255134
rect 548448 254866 548768 254898
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 24114 205774 24734 241218
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 41568 223174 41888 223206
rect 41568 222938 41610 223174
rect 41846 222938 41888 223174
rect 41568 222854 41888 222938
rect 41568 222618 41610 222854
rect 41846 222618 41888 222854
rect 41568 222586 41888 222618
rect 72288 223174 72608 223206
rect 72288 222938 72330 223174
rect 72566 222938 72608 223174
rect 72288 222854 72608 222938
rect 72288 222618 72330 222854
rect 72566 222618 72608 222854
rect 72288 222586 72608 222618
rect 103008 223174 103328 223206
rect 103008 222938 103050 223174
rect 103286 222938 103328 223174
rect 103008 222854 103328 222938
rect 103008 222618 103050 222854
rect 103286 222618 103328 222854
rect 103008 222586 103328 222618
rect 133728 223174 134048 223206
rect 133728 222938 133770 223174
rect 134006 222938 134048 223174
rect 133728 222854 134048 222938
rect 133728 222618 133770 222854
rect 134006 222618 134048 222854
rect 133728 222586 134048 222618
rect 164448 223174 164768 223206
rect 164448 222938 164490 223174
rect 164726 222938 164768 223174
rect 164448 222854 164768 222938
rect 164448 222618 164490 222854
rect 164726 222618 164768 222854
rect 164448 222586 164768 222618
rect 195168 223174 195488 223206
rect 195168 222938 195210 223174
rect 195446 222938 195488 223174
rect 195168 222854 195488 222938
rect 195168 222618 195210 222854
rect 195446 222618 195488 222854
rect 195168 222586 195488 222618
rect 225888 223174 226208 223206
rect 225888 222938 225930 223174
rect 226166 222938 226208 223174
rect 225888 222854 226208 222938
rect 225888 222618 225930 222854
rect 226166 222618 226208 222854
rect 225888 222586 226208 222618
rect 256608 223174 256928 223206
rect 256608 222938 256650 223174
rect 256886 222938 256928 223174
rect 256608 222854 256928 222938
rect 256608 222618 256650 222854
rect 256886 222618 256928 222854
rect 256608 222586 256928 222618
rect 287328 223174 287648 223206
rect 287328 222938 287370 223174
rect 287606 222938 287648 223174
rect 287328 222854 287648 222938
rect 287328 222618 287370 222854
rect 287606 222618 287648 222854
rect 287328 222586 287648 222618
rect 318048 223174 318368 223206
rect 318048 222938 318090 223174
rect 318326 222938 318368 223174
rect 318048 222854 318368 222938
rect 318048 222618 318090 222854
rect 318326 222618 318368 222854
rect 318048 222586 318368 222618
rect 348768 223174 349088 223206
rect 348768 222938 348810 223174
rect 349046 222938 349088 223174
rect 348768 222854 349088 222938
rect 348768 222618 348810 222854
rect 349046 222618 349088 222854
rect 348768 222586 349088 222618
rect 379488 223174 379808 223206
rect 379488 222938 379530 223174
rect 379766 222938 379808 223174
rect 379488 222854 379808 222938
rect 379488 222618 379530 222854
rect 379766 222618 379808 222854
rect 379488 222586 379808 222618
rect 410208 223174 410528 223206
rect 410208 222938 410250 223174
rect 410486 222938 410528 223174
rect 410208 222854 410528 222938
rect 410208 222618 410250 222854
rect 410486 222618 410528 222854
rect 410208 222586 410528 222618
rect 440928 223174 441248 223206
rect 440928 222938 440970 223174
rect 441206 222938 441248 223174
rect 440928 222854 441248 222938
rect 440928 222618 440970 222854
rect 441206 222618 441248 222854
rect 440928 222586 441248 222618
rect 471648 223174 471968 223206
rect 471648 222938 471690 223174
rect 471926 222938 471968 223174
rect 471648 222854 471968 222938
rect 471648 222618 471690 222854
rect 471926 222618 471968 222854
rect 471648 222586 471968 222618
rect 502368 223174 502688 223206
rect 502368 222938 502410 223174
rect 502646 222938 502688 223174
rect 502368 222854 502688 222938
rect 502368 222618 502410 222854
rect 502646 222618 502688 222854
rect 502368 222586 502688 222618
rect 533088 223174 533408 223206
rect 533088 222938 533130 223174
rect 533366 222938 533408 223174
rect 533088 222854 533408 222938
rect 533088 222618 533130 222854
rect 533366 222618 533408 222854
rect 533088 222586 533408 222618
rect 26208 219454 26528 219486
rect 26208 219218 26250 219454
rect 26486 219218 26528 219454
rect 26208 219134 26528 219218
rect 26208 218898 26250 219134
rect 26486 218898 26528 219134
rect 26208 218866 26528 218898
rect 56928 219454 57248 219486
rect 56928 219218 56970 219454
rect 57206 219218 57248 219454
rect 56928 219134 57248 219218
rect 56928 218898 56970 219134
rect 57206 218898 57248 219134
rect 56928 218866 57248 218898
rect 87648 219454 87968 219486
rect 87648 219218 87690 219454
rect 87926 219218 87968 219454
rect 87648 219134 87968 219218
rect 87648 218898 87690 219134
rect 87926 218898 87968 219134
rect 87648 218866 87968 218898
rect 118368 219454 118688 219486
rect 118368 219218 118410 219454
rect 118646 219218 118688 219454
rect 118368 219134 118688 219218
rect 118368 218898 118410 219134
rect 118646 218898 118688 219134
rect 118368 218866 118688 218898
rect 149088 219454 149408 219486
rect 149088 219218 149130 219454
rect 149366 219218 149408 219454
rect 149088 219134 149408 219218
rect 149088 218898 149130 219134
rect 149366 218898 149408 219134
rect 149088 218866 149408 218898
rect 179808 219454 180128 219486
rect 179808 219218 179850 219454
rect 180086 219218 180128 219454
rect 179808 219134 180128 219218
rect 179808 218898 179850 219134
rect 180086 218898 180128 219134
rect 179808 218866 180128 218898
rect 210528 219454 210848 219486
rect 210528 219218 210570 219454
rect 210806 219218 210848 219454
rect 210528 219134 210848 219218
rect 210528 218898 210570 219134
rect 210806 218898 210848 219134
rect 210528 218866 210848 218898
rect 241248 219454 241568 219486
rect 241248 219218 241290 219454
rect 241526 219218 241568 219454
rect 241248 219134 241568 219218
rect 241248 218898 241290 219134
rect 241526 218898 241568 219134
rect 241248 218866 241568 218898
rect 271968 219454 272288 219486
rect 271968 219218 272010 219454
rect 272246 219218 272288 219454
rect 271968 219134 272288 219218
rect 271968 218898 272010 219134
rect 272246 218898 272288 219134
rect 271968 218866 272288 218898
rect 302688 219454 303008 219486
rect 302688 219218 302730 219454
rect 302966 219218 303008 219454
rect 302688 219134 303008 219218
rect 302688 218898 302730 219134
rect 302966 218898 303008 219134
rect 302688 218866 303008 218898
rect 333408 219454 333728 219486
rect 333408 219218 333450 219454
rect 333686 219218 333728 219454
rect 333408 219134 333728 219218
rect 333408 218898 333450 219134
rect 333686 218898 333728 219134
rect 333408 218866 333728 218898
rect 364128 219454 364448 219486
rect 364128 219218 364170 219454
rect 364406 219218 364448 219454
rect 364128 219134 364448 219218
rect 364128 218898 364170 219134
rect 364406 218898 364448 219134
rect 364128 218866 364448 218898
rect 394848 219454 395168 219486
rect 394848 219218 394890 219454
rect 395126 219218 395168 219454
rect 394848 219134 395168 219218
rect 394848 218898 394890 219134
rect 395126 218898 395168 219134
rect 394848 218866 395168 218898
rect 425568 219454 425888 219486
rect 425568 219218 425610 219454
rect 425846 219218 425888 219454
rect 425568 219134 425888 219218
rect 425568 218898 425610 219134
rect 425846 218898 425888 219134
rect 425568 218866 425888 218898
rect 456288 219454 456608 219486
rect 456288 219218 456330 219454
rect 456566 219218 456608 219454
rect 456288 219134 456608 219218
rect 456288 218898 456330 219134
rect 456566 218898 456608 219134
rect 456288 218866 456608 218898
rect 487008 219454 487328 219486
rect 487008 219218 487050 219454
rect 487286 219218 487328 219454
rect 487008 219134 487328 219218
rect 487008 218898 487050 219134
rect 487286 218898 487328 219134
rect 487008 218866 487328 218898
rect 517728 219454 518048 219486
rect 517728 219218 517770 219454
rect 518006 219218 518048 219454
rect 517728 219134 518048 219218
rect 517728 218898 517770 219134
rect 518006 218898 518048 219134
rect 517728 218866 518048 218898
rect 548448 219454 548768 219486
rect 548448 219218 548490 219454
rect 548726 219218 548768 219454
rect 548448 219134 548768 219218
rect 548448 218898 548490 219134
rect 548726 218898 548768 219134
rect 548448 218866 548768 218898
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 24114 169774 24734 205218
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 41568 187174 41888 187206
rect 41568 186938 41610 187174
rect 41846 186938 41888 187174
rect 41568 186854 41888 186938
rect 41568 186618 41610 186854
rect 41846 186618 41888 186854
rect 41568 186586 41888 186618
rect 72288 187174 72608 187206
rect 72288 186938 72330 187174
rect 72566 186938 72608 187174
rect 72288 186854 72608 186938
rect 72288 186618 72330 186854
rect 72566 186618 72608 186854
rect 72288 186586 72608 186618
rect 103008 187174 103328 187206
rect 103008 186938 103050 187174
rect 103286 186938 103328 187174
rect 103008 186854 103328 186938
rect 103008 186618 103050 186854
rect 103286 186618 103328 186854
rect 103008 186586 103328 186618
rect 133728 187174 134048 187206
rect 133728 186938 133770 187174
rect 134006 186938 134048 187174
rect 133728 186854 134048 186938
rect 133728 186618 133770 186854
rect 134006 186618 134048 186854
rect 133728 186586 134048 186618
rect 164448 187174 164768 187206
rect 164448 186938 164490 187174
rect 164726 186938 164768 187174
rect 164448 186854 164768 186938
rect 164448 186618 164490 186854
rect 164726 186618 164768 186854
rect 164448 186586 164768 186618
rect 195168 187174 195488 187206
rect 195168 186938 195210 187174
rect 195446 186938 195488 187174
rect 195168 186854 195488 186938
rect 195168 186618 195210 186854
rect 195446 186618 195488 186854
rect 195168 186586 195488 186618
rect 225888 187174 226208 187206
rect 225888 186938 225930 187174
rect 226166 186938 226208 187174
rect 225888 186854 226208 186938
rect 225888 186618 225930 186854
rect 226166 186618 226208 186854
rect 225888 186586 226208 186618
rect 256608 187174 256928 187206
rect 256608 186938 256650 187174
rect 256886 186938 256928 187174
rect 256608 186854 256928 186938
rect 256608 186618 256650 186854
rect 256886 186618 256928 186854
rect 256608 186586 256928 186618
rect 287328 187174 287648 187206
rect 287328 186938 287370 187174
rect 287606 186938 287648 187174
rect 287328 186854 287648 186938
rect 287328 186618 287370 186854
rect 287606 186618 287648 186854
rect 287328 186586 287648 186618
rect 318048 187174 318368 187206
rect 318048 186938 318090 187174
rect 318326 186938 318368 187174
rect 318048 186854 318368 186938
rect 318048 186618 318090 186854
rect 318326 186618 318368 186854
rect 318048 186586 318368 186618
rect 348768 187174 349088 187206
rect 348768 186938 348810 187174
rect 349046 186938 349088 187174
rect 348768 186854 349088 186938
rect 348768 186618 348810 186854
rect 349046 186618 349088 186854
rect 348768 186586 349088 186618
rect 379488 187174 379808 187206
rect 379488 186938 379530 187174
rect 379766 186938 379808 187174
rect 379488 186854 379808 186938
rect 379488 186618 379530 186854
rect 379766 186618 379808 186854
rect 379488 186586 379808 186618
rect 410208 187174 410528 187206
rect 410208 186938 410250 187174
rect 410486 186938 410528 187174
rect 410208 186854 410528 186938
rect 410208 186618 410250 186854
rect 410486 186618 410528 186854
rect 410208 186586 410528 186618
rect 440928 187174 441248 187206
rect 440928 186938 440970 187174
rect 441206 186938 441248 187174
rect 440928 186854 441248 186938
rect 440928 186618 440970 186854
rect 441206 186618 441248 186854
rect 440928 186586 441248 186618
rect 471648 187174 471968 187206
rect 471648 186938 471690 187174
rect 471926 186938 471968 187174
rect 471648 186854 471968 186938
rect 471648 186618 471690 186854
rect 471926 186618 471968 186854
rect 471648 186586 471968 186618
rect 502368 187174 502688 187206
rect 502368 186938 502410 187174
rect 502646 186938 502688 187174
rect 502368 186854 502688 186938
rect 502368 186618 502410 186854
rect 502646 186618 502688 186854
rect 502368 186586 502688 186618
rect 533088 187174 533408 187206
rect 533088 186938 533130 187174
rect 533366 186938 533408 187174
rect 533088 186854 533408 186938
rect 533088 186618 533130 186854
rect 533366 186618 533408 186854
rect 533088 186586 533408 186618
rect 26208 183454 26528 183486
rect 26208 183218 26250 183454
rect 26486 183218 26528 183454
rect 26208 183134 26528 183218
rect 26208 182898 26250 183134
rect 26486 182898 26528 183134
rect 26208 182866 26528 182898
rect 56928 183454 57248 183486
rect 56928 183218 56970 183454
rect 57206 183218 57248 183454
rect 56928 183134 57248 183218
rect 56928 182898 56970 183134
rect 57206 182898 57248 183134
rect 56928 182866 57248 182898
rect 87648 183454 87968 183486
rect 87648 183218 87690 183454
rect 87926 183218 87968 183454
rect 87648 183134 87968 183218
rect 87648 182898 87690 183134
rect 87926 182898 87968 183134
rect 87648 182866 87968 182898
rect 118368 183454 118688 183486
rect 118368 183218 118410 183454
rect 118646 183218 118688 183454
rect 118368 183134 118688 183218
rect 118368 182898 118410 183134
rect 118646 182898 118688 183134
rect 118368 182866 118688 182898
rect 149088 183454 149408 183486
rect 149088 183218 149130 183454
rect 149366 183218 149408 183454
rect 149088 183134 149408 183218
rect 149088 182898 149130 183134
rect 149366 182898 149408 183134
rect 149088 182866 149408 182898
rect 179808 183454 180128 183486
rect 179808 183218 179850 183454
rect 180086 183218 180128 183454
rect 179808 183134 180128 183218
rect 179808 182898 179850 183134
rect 180086 182898 180128 183134
rect 179808 182866 180128 182898
rect 210528 183454 210848 183486
rect 210528 183218 210570 183454
rect 210806 183218 210848 183454
rect 210528 183134 210848 183218
rect 210528 182898 210570 183134
rect 210806 182898 210848 183134
rect 210528 182866 210848 182898
rect 241248 183454 241568 183486
rect 241248 183218 241290 183454
rect 241526 183218 241568 183454
rect 241248 183134 241568 183218
rect 241248 182898 241290 183134
rect 241526 182898 241568 183134
rect 241248 182866 241568 182898
rect 271968 183454 272288 183486
rect 271968 183218 272010 183454
rect 272246 183218 272288 183454
rect 271968 183134 272288 183218
rect 271968 182898 272010 183134
rect 272246 182898 272288 183134
rect 271968 182866 272288 182898
rect 302688 183454 303008 183486
rect 302688 183218 302730 183454
rect 302966 183218 303008 183454
rect 302688 183134 303008 183218
rect 302688 182898 302730 183134
rect 302966 182898 303008 183134
rect 302688 182866 303008 182898
rect 333408 183454 333728 183486
rect 333408 183218 333450 183454
rect 333686 183218 333728 183454
rect 333408 183134 333728 183218
rect 333408 182898 333450 183134
rect 333686 182898 333728 183134
rect 333408 182866 333728 182898
rect 364128 183454 364448 183486
rect 364128 183218 364170 183454
rect 364406 183218 364448 183454
rect 364128 183134 364448 183218
rect 364128 182898 364170 183134
rect 364406 182898 364448 183134
rect 364128 182866 364448 182898
rect 394848 183454 395168 183486
rect 394848 183218 394890 183454
rect 395126 183218 395168 183454
rect 394848 183134 395168 183218
rect 394848 182898 394890 183134
rect 395126 182898 395168 183134
rect 394848 182866 395168 182898
rect 425568 183454 425888 183486
rect 425568 183218 425610 183454
rect 425846 183218 425888 183454
rect 425568 183134 425888 183218
rect 425568 182898 425610 183134
rect 425846 182898 425888 183134
rect 425568 182866 425888 182898
rect 456288 183454 456608 183486
rect 456288 183218 456330 183454
rect 456566 183218 456608 183454
rect 456288 183134 456608 183218
rect 456288 182898 456330 183134
rect 456566 182898 456608 183134
rect 456288 182866 456608 182898
rect 487008 183454 487328 183486
rect 487008 183218 487050 183454
rect 487286 183218 487328 183454
rect 487008 183134 487328 183218
rect 487008 182898 487050 183134
rect 487286 182898 487328 183134
rect 487008 182866 487328 182898
rect 517728 183454 518048 183486
rect 517728 183218 517770 183454
rect 518006 183218 518048 183454
rect 517728 183134 518048 183218
rect 517728 182898 517770 183134
rect 518006 182898 518048 183134
rect 517728 182866 518048 182898
rect 548448 183454 548768 183486
rect 548448 183218 548490 183454
rect 548726 183218 548768 183454
rect 548448 183134 548768 183218
rect 548448 182898 548490 183134
rect 548726 182898 548768 183134
rect 548448 182866 548768 182898
rect 24114 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 24734 169774
rect 24114 169454 24734 169538
rect 24114 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 24734 169454
rect 24114 133774 24734 169218
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 41568 151174 41888 151206
rect 41568 150938 41610 151174
rect 41846 150938 41888 151174
rect 41568 150854 41888 150938
rect 41568 150618 41610 150854
rect 41846 150618 41888 150854
rect 41568 150586 41888 150618
rect 72288 151174 72608 151206
rect 72288 150938 72330 151174
rect 72566 150938 72608 151174
rect 72288 150854 72608 150938
rect 72288 150618 72330 150854
rect 72566 150618 72608 150854
rect 72288 150586 72608 150618
rect 103008 151174 103328 151206
rect 103008 150938 103050 151174
rect 103286 150938 103328 151174
rect 103008 150854 103328 150938
rect 103008 150618 103050 150854
rect 103286 150618 103328 150854
rect 103008 150586 103328 150618
rect 133728 151174 134048 151206
rect 133728 150938 133770 151174
rect 134006 150938 134048 151174
rect 133728 150854 134048 150938
rect 133728 150618 133770 150854
rect 134006 150618 134048 150854
rect 133728 150586 134048 150618
rect 164448 151174 164768 151206
rect 164448 150938 164490 151174
rect 164726 150938 164768 151174
rect 164448 150854 164768 150938
rect 164448 150618 164490 150854
rect 164726 150618 164768 150854
rect 164448 150586 164768 150618
rect 195168 151174 195488 151206
rect 195168 150938 195210 151174
rect 195446 150938 195488 151174
rect 195168 150854 195488 150938
rect 195168 150618 195210 150854
rect 195446 150618 195488 150854
rect 195168 150586 195488 150618
rect 225888 151174 226208 151206
rect 225888 150938 225930 151174
rect 226166 150938 226208 151174
rect 225888 150854 226208 150938
rect 225888 150618 225930 150854
rect 226166 150618 226208 150854
rect 225888 150586 226208 150618
rect 256608 151174 256928 151206
rect 256608 150938 256650 151174
rect 256886 150938 256928 151174
rect 256608 150854 256928 150938
rect 256608 150618 256650 150854
rect 256886 150618 256928 150854
rect 256608 150586 256928 150618
rect 287328 151174 287648 151206
rect 287328 150938 287370 151174
rect 287606 150938 287648 151174
rect 287328 150854 287648 150938
rect 287328 150618 287370 150854
rect 287606 150618 287648 150854
rect 287328 150586 287648 150618
rect 318048 151174 318368 151206
rect 318048 150938 318090 151174
rect 318326 150938 318368 151174
rect 318048 150854 318368 150938
rect 318048 150618 318090 150854
rect 318326 150618 318368 150854
rect 318048 150586 318368 150618
rect 348768 151174 349088 151206
rect 348768 150938 348810 151174
rect 349046 150938 349088 151174
rect 348768 150854 349088 150938
rect 348768 150618 348810 150854
rect 349046 150618 349088 150854
rect 348768 150586 349088 150618
rect 379488 151174 379808 151206
rect 379488 150938 379530 151174
rect 379766 150938 379808 151174
rect 379488 150854 379808 150938
rect 379488 150618 379530 150854
rect 379766 150618 379808 150854
rect 379488 150586 379808 150618
rect 410208 151174 410528 151206
rect 410208 150938 410250 151174
rect 410486 150938 410528 151174
rect 410208 150854 410528 150938
rect 410208 150618 410250 150854
rect 410486 150618 410528 150854
rect 410208 150586 410528 150618
rect 440928 151174 441248 151206
rect 440928 150938 440970 151174
rect 441206 150938 441248 151174
rect 440928 150854 441248 150938
rect 440928 150618 440970 150854
rect 441206 150618 441248 150854
rect 440928 150586 441248 150618
rect 471648 151174 471968 151206
rect 471648 150938 471690 151174
rect 471926 150938 471968 151174
rect 471648 150854 471968 150938
rect 471648 150618 471690 150854
rect 471926 150618 471968 150854
rect 471648 150586 471968 150618
rect 502368 151174 502688 151206
rect 502368 150938 502410 151174
rect 502646 150938 502688 151174
rect 502368 150854 502688 150938
rect 502368 150618 502410 150854
rect 502646 150618 502688 150854
rect 502368 150586 502688 150618
rect 533088 151174 533408 151206
rect 533088 150938 533130 151174
rect 533366 150938 533408 151174
rect 533088 150854 533408 150938
rect 533088 150618 533130 150854
rect 533366 150618 533408 150854
rect 533088 150586 533408 150618
rect 26208 147454 26528 147486
rect 26208 147218 26250 147454
rect 26486 147218 26528 147454
rect 26208 147134 26528 147218
rect 26208 146898 26250 147134
rect 26486 146898 26528 147134
rect 26208 146866 26528 146898
rect 56928 147454 57248 147486
rect 56928 147218 56970 147454
rect 57206 147218 57248 147454
rect 56928 147134 57248 147218
rect 56928 146898 56970 147134
rect 57206 146898 57248 147134
rect 56928 146866 57248 146898
rect 87648 147454 87968 147486
rect 87648 147218 87690 147454
rect 87926 147218 87968 147454
rect 87648 147134 87968 147218
rect 87648 146898 87690 147134
rect 87926 146898 87968 147134
rect 87648 146866 87968 146898
rect 118368 147454 118688 147486
rect 118368 147218 118410 147454
rect 118646 147218 118688 147454
rect 118368 147134 118688 147218
rect 118368 146898 118410 147134
rect 118646 146898 118688 147134
rect 118368 146866 118688 146898
rect 149088 147454 149408 147486
rect 149088 147218 149130 147454
rect 149366 147218 149408 147454
rect 149088 147134 149408 147218
rect 149088 146898 149130 147134
rect 149366 146898 149408 147134
rect 149088 146866 149408 146898
rect 179808 147454 180128 147486
rect 179808 147218 179850 147454
rect 180086 147218 180128 147454
rect 179808 147134 180128 147218
rect 179808 146898 179850 147134
rect 180086 146898 180128 147134
rect 179808 146866 180128 146898
rect 210528 147454 210848 147486
rect 210528 147218 210570 147454
rect 210806 147218 210848 147454
rect 210528 147134 210848 147218
rect 210528 146898 210570 147134
rect 210806 146898 210848 147134
rect 210528 146866 210848 146898
rect 241248 147454 241568 147486
rect 241248 147218 241290 147454
rect 241526 147218 241568 147454
rect 241248 147134 241568 147218
rect 241248 146898 241290 147134
rect 241526 146898 241568 147134
rect 241248 146866 241568 146898
rect 271968 147454 272288 147486
rect 271968 147218 272010 147454
rect 272246 147218 272288 147454
rect 271968 147134 272288 147218
rect 271968 146898 272010 147134
rect 272246 146898 272288 147134
rect 271968 146866 272288 146898
rect 302688 147454 303008 147486
rect 302688 147218 302730 147454
rect 302966 147218 303008 147454
rect 302688 147134 303008 147218
rect 302688 146898 302730 147134
rect 302966 146898 303008 147134
rect 302688 146866 303008 146898
rect 333408 147454 333728 147486
rect 333408 147218 333450 147454
rect 333686 147218 333728 147454
rect 333408 147134 333728 147218
rect 333408 146898 333450 147134
rect 333686 146898 333728 147134
rect 333408 146866 333728 146898
rect 364128 147454 364448 147486
rect 364128 147218 364170 147454
rect 364406 147218 364448 147454
rect 364128 147134 364448 147218
rect 364128 146898 364170 147134
rect 364406 146898 364448 147134
rect 364128 146866 364448 146898
rect 394848 147454 395168 147486
rect 394848 147218 394890 147454
rect 395126 147218 395168 147454
rect 394848 147134 395168 147218
rect 394848 146898 394890 147134
rect 395126 146898 395168 147134
rect 394848 146866 395168 146898
rect 425568 147454 425888 147486
rect 425568 147218 425610 147454
rect 425846 147218 425888 147454
rect 425568 147134 425888 147218
rect 425568 146898 425610 147134
rect 425846 146898 425888 147134
rect 425568 146866 425888 146898
rect 456288 147454 456608 147486
rect 456288 147218 456330 147454
rect 456566 147218 456608 147454
rect 456288 147134 456608 147218
rect 456288 146898 456330 147134
rect 456566 146898 456608 147134
rect 456288 146866 456608 146898
rect 487008 147454 487328 147486
rect 487008 147218 487050 147454
rect 487286 147218 487328 147454
rect 487008 147134 487328 147218
rect 487008 146898 487050 147134
rect 487286 146898 487328 147134
rect 487008 146866 487328 146898
rect 517728 147454 518048 147486
rect 517728 147218 517770 147454
rect 518006 147218 518048 147454
rect 517728 147134 518048 147218
rect 517728 146898 517770 147134
rect 518006 146898 518048 147134
rect 517728 146866 518048 146898
rect 548448 147454 548768 147486
rect 548448 147218 548490 147454
rect 548726 147218 548768 147454
rect 548448 147134 548768 147218
rect 548448 146898 548490 147134
rect 548726 146898 548768 147134
rect 548448 146866 548768 146898
rect 24114 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 24734 133774
rect 24114 133454 24734 133538
rect 24114 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 24734 133454
rect 24114 97774 24734 133218
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 41568 115174 41888 115206
rect 41568 114938 41610 115174
rect 41846 114938 41888 115174
rect 41568 114854 41888 114938
rect 41568 114618 41610 114854
rect 41846 114618 41888 114854
rect 41568 114586 41888 114618
rect 72288 115174 72608 115206
rect 72288 114938 72330 115174
rect 72566 114938 72608 115174
rect 72288 114854 72608 114938
rect 72288 114618 72330 114854
rect 72566 114618 72608 114854
rect 72288 114586 72608 114618
rect 103008 115174 103328 115206
rect 103008 114938 103050 115174
rect 103286 114938 103328 115174
rect 103008 114854 103328 114938
rect 103008 114618 103050 114854
rect 103286 114618 103328 114854
rect 103008 114586 103328 114618
rect 133728 115174 134048 115206
rect 133728 114938 133770 115174
rect 134006 114938 134048 115174
rect 133728 114854 134048 114938
rect 133728 114618 133770 114854
rect 134006 114618 134048 114854
rect 133728 114586 134048 114618
rect 164448 115174 164768 115206
rect 164448 114938 164490 115174
rect 164726 114938 164768 115174
rect 164448 114854 164768 114938
rect 164448 114618 164490 114854
rect 164726 114618 164768 114854
rect 164448 114586 164768 114618
rect 195168 115174 195488 115206
rect 195168 114938 195210 115174
rect 195446 114938 195488 115174
rect 195168 114854 195488 114938
rect 195168 114618 195210 114854
rect 195446 114618 195488 114854
rect 195168 114586 195488 114618
rect 225888 115174 226208 115206
rect 225888 114938 225930 115174
rect 226166 114938 226208 115174
rect 225888 114854 226208 114938
rect 225888 114618 225930 114854
rect 226166 114618 226208 114854
rect 225888 114586 226208 114618
rect 256608 115174 256928 115206
rect 256608 114938 256650 115174
rect 256886 114938 256928 115174
rect 256608 114854 256928 114938
rect 256608 114618 256650 114854
rect 256886 114618 256928 114854
rect 256608 114586 256928 114618
rect 287328 115174 287648 115206
rect 287328 114938 287370 115174
rect 287606 114938 287648 115174
rect 287328 114854 287648 114938
rect 287328 114618 287370 114854
rect 287606 114618 287648 114854
rect 287328 114586 287648 114618
rect 318048 115174 318368 115206
rect 318048 114938 318090 115174
rect 318326 114938 318368 115174
rect 318048 114854 318368 114938
rect 318048 114618 318090 114854
rect 318326 114618 318368 114854
rect 318048 114586 318368 114618
rect 348768 115174 349088 115206
rect 348768 114938 348810 115174
rect 349046 114938 349088 115174
rect 348768 114854 349088 114938
rect 348768 114618 348810 114854
rect 349046 114618 349088 114854
rect 348768 114586 349088 114618
rect 379488 115174 379808 115206
rect 379488 114938 379530 115174
rect 379766 114938 379808 115174
rect 379488 114854 379808 114938
rect 379488 114618 379530 114854
rect 379766 114618 379808 114854
rect 379488 114586 379808 114618
rect 410208 115174 410528 115206
rect 410208 114938 410250 115174
rect 410486 114938 410528 115174
rect 410208 114854 410528 114938
rect 410208 114618 410250 114854
rect 410486 114618 410528 114854
rect 410208 114586 410528 114618
rect 440928 115174 441248 115206
rect 440928 114938 440970 115174
rect 441206 114938 441248 115174
rect 440928 114854 441248 114938
rect 440928 114618 440970 114854
rect 441206 114618 441248 114854
rect 440928 114586 441248 114618
rect 471648 115174 471968 115206
rect 471648 114938 471690 115174
rect 471926 114938 471968 115174
rect 471648 114854 471968 114938
rect 471648 114618 471690 114854
rect 471926 114618 471968 114854
rect 471648 114586 471968 114618
rect 502368 115174 502688 115206
rect 502368 114938 502410 115174
rect 502646 114938 502688 115174
rect 502368 114854 502688 114938
rect 502368 114618 502410 114854
rect 502646 114618 502688 114854
rect 502368 114586 502688 114618
rect 533088 115174 533408 115206
rect 533088 114938 533130 115174
rect 533366 114938 533408 115174
rect 533088 114854 533408 114938
rect 533088 114618 533130 114854
rect 533366 114618 533408 114854
rect 533088 114586 533408 114618
rect 26208 111454 26528 111486
rect 26208 111218 26250 111454
rect 26486 111218 26528 111454
rect 26208 111134 26528 111218
rect 26208 110898 26250 111134
rect 26486 110898 26528 111134
rect 26208 110866 26528 110898
rect 56928 111454 57248 111486
rect 56928 111218 56970 111454
rect 57206 111218 57248 111454
rect 56928 111134 57248 111218
rect 56928 110898 56970 111134
rect 57206 110898 57248 111134
rect 56928 110866 57248 110898
rect 87648 111454 87968 111486
rect 87648 111218 87690 111454
rect 87926 111218 87968 111454
rect 87648 111134 87968 111218
rect 87648 110898 87690 111134
rect 87926 110898 87968 111134
rect 87648 110866 87968 110898
rect 118368 111454 118688 111486
rect 118368 111218 118410 111454
rect 118646 111218 118688 111454
rect 118368 111134 118688 111218
rect 118368 110898 118410 111134
rect 118646 110898 118688 111134
rect 118368 110866 118688 110898
rect 149088 111454 149408 111486
rect 149088 111218 149130 111454
rect 149366 111218 149408 111454
rect 149088 111134 149408 111218
rect 149088 110898 149130 111134
rect 149366 110898 149408 111134
rect 149088 110866 149408 110898
rect 179808 111454 180128 111486
rect 179808 111218 179850 111454
rect 180086 111218 180128 111454
rect 179808 111134 180128 111218
rect 179808 110898 179850 111134
rect 180086 110898 180128 111134
rect 179808 110866 180128 110898
rect 210528 111454 210848 111486
rect 210528 111218 210570 111454
rect 210806 111218 210848 111454
rect 210528 111134 210848 111218
rect 210528 110898 210570 111134
rect 210806 110898 210848 111134
rect 210528 110866 210848 110898
rect 241248 111454 241568 111486
rect 241248 111218 241290 111454
rect 241526 111218 241568 111454
rect 241248 111134 241568 111218
rect 241248 110898 241290 111134
rect 241526 110898 241568 111134
rect 241248 110866 241568 110898
rect 271968 111454 272288 111486
rect 271968 111218 272010 111454
rect 272246 111218 272288 111454
rect 271968 111134 272288 111218
rect 271968 110898 272010 111134
rect 272246 110898 272288 111134
rect 271968 110866 272288 110898
rect 302688 111454 303008 111486
rect 302688 111218 302730 111454
rect 302966 111218 303008 111454
rect 302688 111134 303008 111218
rect 302688 110898 302730 111134
rect 302966 110898 303008 111134
rect 302688 110866 303008 110898
rect 333408 111454 333728 111486
rect 333408 111218 333450 111454
rect 333686 111218 333728 111454
rect 333408 111134 333728 111218
rect 333408 110898 333450 111134
rect 333686 110898 333728 111134
rect 333408 110866 333728 110898
rect 364128 111454 364448 111486
rect 364128 111218 364170 111454
rect 364406 111218 364448 111454
rect 364128 111134 364448 111218
rect 364128 110898 364170 111134
rect 364406 110898 364448 111134
rect 364128 110866 364448 110898
rect 394848 111454 395168 111486
rect 394848 111218 394890 111454
rect 395126 111218 395168 111454
rect 394848 111134 395168 111218
rect 394848 110898 394890 111134
rect 395126 110898 395168 111134
rect 394848 110866 395168 110898
rect 425568 111454 425888 111486
rect 425568 111218 425610 111454
rect 425846 111218 425888 111454
rect 425568 111134 425888 111218
rect 425568 110898 425610 111134
rect 425846 110898 425888 111134
rect 425568 110866 425888 110898
rect 456288 111454 456608 111486
rect 456288 111218 456330 111454
rect 456566 111218 456608 111454
rect 456288 111134 456608 111218
rect 456288 110898 456330 111134
rect 456566 110898 456608 111134
rect 456288 110866 456608 110898
rect 487008 111454 487328 111486
rect 487008 111218 487050 111454
rect 487286 111218 487328 111454
rect 487008 111134 487328 111218
rect 487008 110898 487050 111134
rect 487286 110898 487328 111134
rect 487008 110866 487328 110898
rect 517728 111454 518048 111486
rect 517728 111218 517770 111454
rect 518006 111218 518048 111454
rect 517728 111134 518048 111218
rect 517728 110898 517770 111134
rect 518006 110898 518048 111134
rect 517728 110866 518048 110898
rect 548448 111454 548768 111486
rect 548448 111218 548490 111454
rect 548726 111218 548768 111454
rect 548448 111134 548768 111218
rect 548448 110898 548490 111134
rect 548726 110898 548768 111134
rect 548448 110866 548768 110898
rect 24114 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 24734 97774
rect 24114 97454 24734 97538
rect 24114 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 24734 97454
rect 24114 61774 24734 97218
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 41568 79174 41888 79206
rect 41568 78938 41610 79174
rect 41846 78938 41888 79174
rect 41568 78854 41888 78938
rect 41568 78618 41610 78854
rect 41846 78618 41888 78854
rect 41568 78586 41888 78618
rect 72288 79174 72608 79206
rect 72288 78938 72330 79174
rect 72566 78938 72608 79174
rect 72288 78854 72608 78938
rect 72288 78618 72330 78854
rect 72566 78618 72608 78854
rect 72288 78586 72608 78618
rect 103008 79174 103328 79206
rect 103008 78938 103050 79174
rect 103286 78938 103328 79174
rect 103008 78854 103328 78938
rect 103008 78618 103050 78854
rect 103286 78618 103328 78854
rect 103008 78586 103328 78618
rect 133728 79174 134048 79206
rect 133728 78938 133770 79174
rect 134006 78938 134048 79174
rect 133728 78854 134048 78938
rect 133728 78618 133770 78854
rect 134006 78618 134048 78854
rect 133728 78586 134048 78618
rect 164448 79174 164768 79206
rect 164448 78938 164490 79174
rect 164726 78938 164768 79174
rect 164448 78854 164768 78938
rect 164448 78618 164490 78854
rect 164726 78618 164768 78854
rect 164448 78586 164768 78618
rect 195168 79174 195488 79206
rect 195168 78938 195210 79174
rect 195446 78938 195488 79174
rect 195168 78854 195488 78938
rect 195168 78618 195210 78854
rect 195446 78618 195488 78854
rect 195168 78586 195488 78618
rect 225888 79174 226208 79206
rect 225888 78938 225930 79174
rect 226166 78938 226208 79174
rect 225888 78854 226208 78938
rect 225888 78618 225930 78854
rect 226166 78618 226208 78854
rect 225888 78586 226208 78618
rect 256608 79174 256928 79206
rect 256608 78938 256650 79174
rect 256886 78938 256928 79174
rect 256608 78854 256928 78938
rect 256608 78618 256650 78854
rect 256886 78618 256928 78854
rect 256608 78586 256928 78618
rect 287328 79174 287648 79206
rect 287328 78938 287370 79174
rect 287606 78938 287648 79174
rect 287328 78854 287648 78938
rect 287328 78618 287370 78854
rect 287606 78618 287648 78854
rect 287328 78586 287648 78618
rect 318048 79174 318368 79206
rect 318048 78938 318090 79174
rect 318326 78938 318368 79174
rect 318048 78854 318368 78938
rect 318048 78618 318090 78854
rect 318326 78618 318368 78854
rect 318048 78586 318368 78618
rect 348768 79174 349088 79206
rect 348768 78938 348810 79174
rect 349046 78938 349088 79174
rect 348768 78854 349088 78938
rect 348768 78618 348810 78854
rect 349046 78618 349088 78854
rect 348768 78586 349088 78618
rect 379488 79174 379808 79206
rect 379488 78938 379530 79174
rect 379766 78938 379808 79174
rect 379488 78854 379808 78938
rect 379488 78618 379530 78854
rect 379766 78618 379808 78854
rect 379488 78586 379808 78618
rect 410208 79174 410528 79206
rect 410208 78938 410250 79174
rect 410486 78938 410528 79174
rect 410208 78854 410528 78938
rect 410208 78618 410250 78854
rect 410486 78618 410528 78854
rect 410208 78586 410528 78618
rect 440928 79174 441248 79206
rect 440928 78938 440970 79174
rect 441206 78938 441248 79174
rect 440928 78854 441248 78938
rect 440928 78618 440970 78854
rect 441206 78618 441248 78854
rect 440928 78586 441248 78618
rect 471648 79174 471968 79206
rect 471648 78938 471690 79174
rect 471926 78938 471968 79174
rect 471648 78854 471968 78938
rect 471648 78618 471690 78854
rect 471926 78618 471968 78854
rect 471648 78586 471968 78618
rect 502368 79174 502688 79206
rect 502368 78938 502410 79174
rect 502646 78938 502688 79174
rect 502368 78854 502688 78938
rect 502368 78618 502410 78854
rect 502646 78618 502688 78854
rect 502368 78586 502688 78618
rect 533088 79174 533408 79206
rect 533088 78938 533130 79174
rect 533366 78938 533408 79174
rect 533088 78854 533408 78938
rect 533088 78618 533130 78854
rect 533366 78618 533408 78854
rect 533088 78586 533408 78618
rect 26208 75454 26528 75486
rect 26208 75218 26250 75454
rect 26486 75218 26528 75454
rect 26208 75134 26528 75218
rect 26208 74898 26250 75134
rect 26486 74898 26528 75134
rect 26208 74866 26528 74898
rect 56928 75454 57248 75486
rect 56928 75218 56970 75454
rect 57206 75218 57248 75454
rect 56928 75134 57248 75218
rect 56928 74898 56970 75134
rect 57206 74898 57248 75134
rect 56928 74866 57248 74898
rect 87648 75454 87968 75486
rect 87648 75218 87690 75454
rect 87926 75218 87968 75454
rect 87648 75134 87968 75218
rect 87648 74898 87690 75134
rect 87926 74898 87968 75134
rect 87648 74866 87968 74898
rect 118368 75454 118688 75486
rect 118368 75218 118410 75454
rect 118646 75218 118688 75454
rect 118368 75134 118688 75218
rect 118368 74898 118410 75134
rect 118646 74898 118688 75134
rect 118368 74866 118688 74898
rect 149088 75454 149408 75486
rect 149088 75218 149130 75454
rect 149366 75218 149408 75454
rect 149088 75134 149408 75218
rect 149088 74898 149130 75134
rect 149366 74898 149408 75134
rect 149088 74866 149408 74898
rect 179808 75454 180128 75486
rect 179808 75218 179850 75454
rect 180086 75218 180128 75454
rect 179808 75134 180128 75218
rect 179808 74898 179850 75134
rect 180086 74898 180128 75134
rect 179808 74866 180128 74898
rect 210528 75454 210848 75486
rect 210528 75218 210570 75454
rect 210806 75218 210848 75454
rect 210528 75134 210848 75218
rect 210528 74898 210570 75134
rect 210806 74898 210848 75134
rect 210528 74866 210848 74898
rect 241248 75454 241568 75486
rect 241248 75218 241290 75454
rect 241526 75218 241568 75454
rect 241248 75134 241568 75218
rect 241248 74898 241290 75134
rect 241526 74898 241568 75134
rect 241248 74866 241568 74898
rect 271968 75454 272288 75486
rect 271968 75218 272010 75454
rect 272246 75218 272288 75454
rect 271968 75134 272288 75218
rect 271968 74898 272010 75134
rect 272246 74898 272288 75134
rect 271968 74866 272288 74898
rect 302688 75454 303008 75486
rect 302688 75218 302730 75454
rect 302966 75218 303008 75454
rect 302688 75134 303008 75218
rect 302688 74898 302730 75134
rect 302966 74898 303008 75134
rect 302688 74866 303008 74898
rect 333408 75454 333728 75486
rect 333408 75218 333450 75454
rect 333686 75218 333728 75454
rect 333408 75134 333728 75218
rect 333408 74898 333450 75134
rect 333686 74898 333728 75134
rect 333408 74866 333728 74898
rect 364128 75454 364448 75486
rect 364128 75218 364170 75454
rect 364406 75218 364448 75454
rect 364128 75134 364448 75218
rect 364128 74898 364170 75134
rect 364406 74898 364448 75134
rect 364128 74866 364448 74898
rect 394848 75454 395168 75486
rect 394848 75218 394890 75454
rect 395126 75218 395168 75454
rect 394848 75134 395168 75218
rect 394848 74898 394890 75134
rect 395126 74898 395168 75134
rect 394848 74866 395168 74898
rect 425568 75454 425888 75486
rect 425568 75218 425610 75454
rect 425846 75218 425888 75454
rect 425568 75134 425888 75218
rect 425568 74898 425610 75134
rect 425846 74898 425888 75134
rect 425568 74866 425888 74898
rect 456288 75454 456608 75486
rect 456288 75218 456330 75454
rect 456566 75218 456608 75454
rect 456288 75134 456608 75218
rect 456288 74898 456330 75134
rect 456566 74898 456608 75134
rect 456288 74866 456608 74898
rect 487008 75454 487328 75486
rect 487008 75218 487050 75454
rect 487286 75218 487328 75454
rect 487008 75134 487328 75218
rect 487008 74898 487050 75134
rect 487286 74898 487328 75134
rect 487008 74866 487328 74898
rect 517728 75454 518048 75486
rect 517728 75218 517770 75454
rect 518006 75218 518048 75454
rect 517728 75134 518048 75218
rect 517728 74898 517770 75134
rect 518006 74898 518048 75134
rect 517728 74866 518048 74898
rect 548448 75454 548768 75486
rect 548448 75218 548490 75454
rect 548726 75218 548768 75454
rect 548448 75134 548768 75218
rect 548448 74898 548490 75134
rect 548726 74898 548768 75134
rect 548448 74866 548768 74898
rect 24114 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 24734 61774
rect 24114 61454 24734 61538
rect 24114 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 24734 61454
rect 22507 42940 22573 42941
rect 22507 42876 22508 42940
rect 22572 42876 22573 42940
rect 22507 42875 22573 42876
rect 22510 35910 22570 42875
rect 22510 35850 22754 35910
rect 21955 22676 22021 22677
rect 21955 22612 21956 22676
rect 22020 22612 22021 22676
rect 21955 22611 22021 22612
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20115 5132 20181 5133
rect 20115 5068 20116 5132
rect 20180 5068 20181 5132
rect 20115 5067 20181 5068
rect 19931 4996 19997 4997
rect 19931 4932 19932 4996
rect 19996 4932 19997 4996
rect 19931 4931 19997 4932
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 -5146 21014 21498
rect 22694 21317 22754 35850
rect 24114 25774 24734 61218
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 41568 43174 41888 43206
rect 41568 42938 41610 43174
rect 41846 42938 41888 43174
rect 41568 42854 41888 42938
rect 41568 42618 41610 42854
rect 41846 42618 41888 42854
rect 41568 42586 41888 42618
rect 72288 43174 72608 43206
rect 72288 42938 72330 43174
rect 72566 42938 72608 43174
rect 72288 42854 72608 42938
rect 72288 42618 72330 42854
rect 72566 42618 72608 42854
rect 72288 42586 72608 42618
rect 103008 43174 103328 43206
rect 103008 42938 103050 43174
rect 103286 42938 103328 43174
rect 103008 42854 103328 42938
rect 103008 42618 103050 42854
rect 103286 42618 103328 42854
rect 103008 42586 103328 42618
rect 133728 43174 134048 43206
rect 133728 42938 133770 43174
rect 134006 42938 134048 43174
rect 133728 42854 134048 42938
rect 133728 42618 133770 42854
rect 134006 42618 134048 42854
rect 133728 42586 134048 42618
rect 164448 43174 164768 43206
rect 164448 42938 164490 43174
rect 164726 42938 164768 43174
rect 164448 42854 164768 42938
rect 164448 42618 164490 42854
rect 164726 42618 164768 42854
rect 164448 42586 164768 42618
rect 195168 43174 195488 43206
rect 195168 42938 195210 43174
rect 195446 42938 195488 43174
rect 195168 42854 195488 42938
rect 195168 42618 195210 42854
rect 195446 42618 195488 42854
rect 195168 42586 195488 42618
rect 225888 43174 226208 43206
rect 225888 42938 225930 43174
rect 226166 42938 226208 43174
rect 225888 42854 226208 42938
rect 225888 42618 225930 42854
rect 226166 42618 226208 42854
rect 225888 42586 226208 42618
rect 256608 43174 256928 43206
rect 256608 42938 256650 43174
rect 256886 42938 256928 43174
rect 256608 42854 256928 42938
rect 256608 42618 256650 42854
rect 256886 42618 256928 42854
rect 256608 42586 256928 42618
rect 287328 43174 287648 43206
rect 287328 42938 287370 43174
rect 287606 42938 287648 43174
rect 287328 42854 287648 42938
rect 287328 42618 287370 42854
rect 287606 42618 287648 42854
rect 287328 42586 287648 42618
rect 318048 43174 318368 43206
rect 318048 42938 318090 43174
rect 318326 42938 318368 43174
rect 318048 42854 318368 42938
rect 318048 42618 318090 42854
rect 318326 42618 318368 42854
rect 318048 42586 318368 42618
rect 348768 43174 349088 43206
rect 348768 42938 348810 43174
rect 349046 42938 349088 43174
rect 348768 42854 349088 42938
rect 348768 42618 348810 42854
rect 349046 42618 349088 42854
rect 348768 42586 349088 42618
rect 379488 43174 379808 43206
rect 379488 42938 379530 43174
rect 379766 42938 379808 43174
rect 379488 42854 379808 42938
rect 379488 42618 379530 42854
rect 379766 42618 379808 42854
rect 379488 42586 379808 42618
rect 410208 43174 410528 43206
rect 410208 42938 410250 43174
rect 410486 42938 410528 43174
rect 410208 42854 410528 42938
rect 410208 42618 410250 42854
rect 410486 42618 410528 42854
rect 410208 42586 410528 42618
rect 440928 43174 441248 43206
rect 440928 42938 440970 43174
rect 441206 42938 441248 43174
rect 440928 42854 441248 42938
rect 440928 42618 440970 42854
rect 441206 42618 441248 42854
rect 440928 42586 441248 42618
rect 471648 43174 471968 43206
rect 471648 42938 471690 43174
rect 471926 42938 471968 43174
rect 471648 42854 471968 42938
rect 471648 42618 471690 42854
rect 471926 42618 471968 42854
rect 471648 42586 471968 42618
rect 502368 43174 502688 43206
rect 502368 42938 502410 43174
rect 502646 42938 502688 43174
rect 502368 42854 502688 42938
rect 502368 42618 502410 42854
rect 502646 42618 502688 42854
rect 502368 42586 502688 42618
rect 533088 43174 533408 43206
rect 533088 42938 533130 43174
rect 533366 42938 533408 43174
rect 533088 42854 533408 42938
rect 533088 42618 533130 42854
rect 533366 42618 533408 42854
rect 533088 42586 533408 42618
rect 26208 39454 26528 39486
rect 26208 39218 26250 39454
rect 26486 39218 26528 39454
rect 26208 39134 26528 39218
rect 26208 38898 26250 39134
rect 26486 38898 26528 39134
rect 26208 38866 26528 38898
rect 56928 39454 57248 39486
rect 56928 39218 56970 39454
rect 57206 39218 57248 39454
rect 56928 39134 57248 39218
rect 56928 38898 56970 39134
rect 57206 38898 57248 39134
rect 56928 38866 57248 38898
rect 87648 39454 87968 39486
rect 87648 39218 87690 39454
rect 87926 39218 87968 39454
rect 87648 39134 87968 39218
rect 87648 38898 87690 39134
rect 87926 38898 87968 39134
rect 87648 38866 87968 38898
rect 118368 39454 118688 39486
rect 118368 39218 118410 39454
rect 118646 39218 118688 39454
rect 118368 39134 118688 39218
rect 118368 38898 118410 39134
rect 118646 38898 118688 39134
rect 118368 38866 118688 38898
rect 149088 39454 149408 39486
rect 149088 39218 149130 39454
rect 149366 39218 149408 39454
rect 149088 39134 149408 39218
rect 149088 38898 149130 39134
rect 149366 38898 149408 39134
rect 149088 38866 149408 38898
rect 179808 39454 180128 39486
rect 179808 39218 179850 39454
rect 180086 39218 180128 39454
rect 179808 39134 180128 39218
rect 179808 38898 179850 39134
rect 180086 38898 180128 39134
rect 179808 38866 180128 38898
rect 210528 39454 210848 39486
rect 210528 39218 210570 39454
rect 210806 39218 210848 39454
rect 210528 39134 210848 39218
rect 210528 38898 210570 39134
rect 210806 38898 210848 39134
rect 210528 38866 210848 38898
rect 241248 39454 241568 39486
rect 241248 39218 241290 39454
rect 241526 39218 241568 39454
rect 241248 39134 241568 39218
rect 241248 38898 241290 39134
rect 241526 38898 241568 39134
rect 241248 38866 241568 38898
rect 271968 39454 272288 39486
rect 271968 39218 272010 39454
rect 272246 39218 272288 39454
rect 271968 39134 272288 39218
rect 271968 38898 272010 39134
rect 272246 38898 272288 39134
rect 271968 38866 272288 38898
rect 302688 39454 303008 39486
rect 302688 39218 302730 39454
rect 302966 39218 303008 39454
rect 302688 39134 303008 39218
rect 302688 38898 302730 39134
rect 302966 38898 303008 39134
rect 302688 38866 303008 38898
rect 333408 39454 333728 39486
rect 333408 39218 333450 39454
rect 333686 39218 333728 39454
rect 333408 39134 333728 39218
rect 333408 38898 333450 39134
rect 333686 38898 333728 39134
rect 333408 38866 333728 38898
rect 364128 39454 364448 39486
rect 364128 39218 364170 39454
rect 364406 39218 364448 39454
rect 364128 39134 364448 39218
rect 364128 38898 364170 39134
rect 364406 38898 364448 39134
rect 364128 38866 364448 38898
rect 394848 39454 395168 39486
rect 394848 39218 394890 39454
rect 395126 39218 395168 39454
rect 394848 39134 395168 39218
rect 394848 38898 394890 39134
rect 395126 38898 395168 39134
rect 394848 38866 395168 38898
rect 425568 39454 425888 39486
rect 425568 39218 425610 39454
rect 425846 39218 425888 39454
rect 425568 39134 425888 39218
rect 425568 38898 425610 39134
rect 425846 38898 425888 39134
rect 425568 38866 425888 38898
rect 456288 39454 456608 39486
rect 456288 39218 456330 39454
rect 456566 39218 456608 39454
rect 456288 39134 456608 39218
rect 456288 38898 456330 39134
rect 456566 38898 456608 39134
rect 456288 38866 456608 38898
rect 487008 39454 487328 39486
rect 487008 39218 487050 39454
rect 487286 39218 487328 39454
rect 487008 39134 487328 39218
rect 487008 38898 487050 39134
rect 487286 38898 487328 39134
rect 487008 38866 487328 38898
rect 517728 39454 518048 39486
rect 517728 39218 517770 39454
rect 518006 39218 518048 39454
rect 517728 39134 518048 39218
rect 517728 38898 517770 39134
rect 518006 38898 518048 39134
rect 517728 38866 518048 38898
rect 548448 39454 548768 39486
rect 548448 39218 548490 39454
rect 548726 39218 548768 39454
rect 548448 39134 548768 39218
rect 548448 38898 548490 39134
rect 548726 38898 548768 39134
rect 548448 38866 548768 38898
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 23795 23492 23861 23493
rect 23795 23428 23796 23492
rect 23860 23428 23861 23492
rect 23795 23427 23861 23428
rect 22691 21316 22757 21317
rect 22691 21252 22692 21316
rect 22756 21252 22757 21316
rect 22691 21251 22757 21252
rect 23798 4045 23858 23427
rect 23795 4044 23861 4045
rect 23795 3980 23796 4044
rect 23860 3980 23861 4044
rect 23795 3979 23861 3980
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 37794 3454 38414 22287
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 7174 42134 22068
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 10894 45854 22287
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 22287
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 18334 53294 22287
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 21885 57014 22068
rect 56394 21649 56426 21885
rect 56662 21649 56746 21885
rect 56982 21649 57014 21885
rect 56394 -5146 57014 21649
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 73794 3454 74414 22287
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 7174 78134 22287
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 10894 81854 22287
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 14614 85574 22287
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 18334 89294 22287
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 22054 93014 22287
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 109794 3454 110414 22287
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 7174 114134 22287
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 10894 117854 22287
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 14614 121574 22287
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 18334 125294 22287
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 22054 129014 22287
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 145794 3454 146414 22287
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 7174 150134 22287
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 10894 153854 22287
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 14614 157574 22287
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 18334 161294 22287
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 21885 165014 22068
rect 164394 21649 164426 21885
rect 164662 21649 164746 21885
rect 164982 21649 165014 21885
rect 164394 -5146 165014 21649
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 181794 3454 182414 22287
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 7174 186134 22287
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 10894 189854 22287
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 22287
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 22287
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 22054 201014 22287
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 217794 3454 218414 22287
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 7174 222134 22287
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 10894 225854 22068
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 14614 229574 22287
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 22287
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 22054 237014 22287
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 253794 3454 254414 22287
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 7174 258134 22287
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 10894 261854 22287
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 14614 265574 22287
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 18334 269294 22287
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 22054 273014 22287
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 289794 3454 290414 22287
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 7174 294134 22287
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 10894 297854 22287
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 22287
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 18334 305294 22287
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 22054 309014 22287
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 325794 3454 326414 22287
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 7174 330134 22287
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 10894 333854 22068
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 14614 337574 22287
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 18334 341294 22287
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 22054 345014 22287
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 361794 3454 362414 22287
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 7174 366134 22287
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 10894 369854 22287
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 14614 373574 22287
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 18334 377294 22287
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 22054 381014 22287
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 397794 3454 398414 22287
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 7174 402134 22287
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 10894 405854 22287
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 14614 409574 22287
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 18334 413294 22287
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 22287
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 433794 3454 434414 22287
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 22287
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 10894 441854 22068
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 14614 445574 22287
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 22287
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 22054 453014 22287
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 469794 3454 470414 22287
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 7174 474134 22287
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 10894 477854 22287
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 14614 481574 22287
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 18334 485294 22287
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 22054 489014 22287
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 505794 3454 506414 22287
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 7174 510134 22287
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 10894 513854 22287
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 14614 517574 22287
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 18334 521294 22287
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 22054 525014 22287
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 541794 3454 542414 22287
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 22287
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 22287
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 22287
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18334 557294 22287
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 561630 4997 561690 659227
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 561811 636172 561877 636173
rect 561811 636108 561812 636172
rect 561876 636108 561877 636172
rect 561811 636107 561877 636108
rect 561627 4996 561693 4997
rect 561627 4932 561628 4996
rect 561692 4932 561693 4996
rect 561627 4931 561693 4932
rect 561814 3773 561874 636107
rect 563099 613732 563165 613733
rect 563099 613668 563100 613732
rect 563164 613668 563165 613732
rect 563099 613667 563165 613668
rect 561995 590068 562061 590069
rect 561995 590004 561996 590068
rect 562060 590004 562061 590068
rect 561995 590003 562061 590004
rect 561998 4861 562058 590003
rect 562179 545052 562245 545053
rect 562179 544988 562180 545052
rect 562244 544988 562245 545052
rect 562179 544987 562245 544988
rect 562182 6357 562242 544987
rect 562179 6356 562245 6357
rect 562179 6292 562180 6356
rect 562244 6292 562245 6356
rect 562179 6291 562245 6292
rect 563102 6221 563162 613667
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 563283 522612 563349 522613
rect 563283 522548 563284 522612
rect 563348 522548 563349 522612
rect 563283 522547 563349 522548
rect 563099 6220 563165 6221
rect 563099 6156 563100 6220
rect 563164 6156 563165 6220
rect 563099 6155 563165 6156
rect 561995 4860 562061 4861
rect 561995 4796 561996 4860
rect 562060 4796 562061 4860
rect 561995 4795 562061 4796
rect 561811 3772 561877 3773
rect 561811 3708 561812 3772
rect 561876 3708 561877 3772
rect 561811 3707 561877 3708
rect 563286 3637 563346 522547
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 563467 453932 563533 453933
rect 563467 453868 563468 453932
rect 563532 453868 563533 453932
rect 563467 453867 563533 453868
rect 563283 3636 563349 3637
rect 563283 3572 563284 3636
rect 563348 3572 563349 3636
rect 563283 3571 563349 3572
rect 563470 3501 563530 453867
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 563467 3500 563533 3501
rect 563467 3436 563468 3500
rect 563532 3436 563533 3500
rect 563467 3435 563533 3436
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 41610 654938 41846 655174
rect 41610 654618 41846 654854
rect 72330 654938 72566 655174
rect 72330 654618 72566 654854
rect 103050 654938 103286 655174
rect 103050 654618 103286 654854
rect 133770 654938 134006 655174
rect 133770 654618 134006 654854
rect 164490 654938 164726 655174
rect 164490 654618 164726 654854
rect 195210 654938 195446 655174
rect 195210 654618 195446 654854
rect 225930 654938 226166 655174
rect 225930 654618 226166 654854
rect 256650 654938 256886 655174
rect 256650 654618 256886 654854
rect 287370 654938 287606 655174
rect 287370 654618 287606 654854
rect 318090 654938 318326 655174
rect 318090 654618 318326 654854
rect 348810 654938 349046 655174
rect 348810 654618 349046 654854
rect 379530 654938 379766 655174
rect 379530 654618 379766 654854
rect 410250 654938 410486 655174
rect 410250 654618 410486 654854
rect 440970 654938 441206 655174
rect 440970 654618 441206 654854
rect 471690 654938 471926 655174
rect 471690 654618 471926 654854
rect 502410 654938 502646 655174
rect 502410 654618 502646 654854
rect 533130 654938 533366 655174
rect 533130 654618 533366 654854
rect 26250 651218 26486 651454
rect 26250 650898 26486 651134
rect 56970 651218 57206 651454
rect 56970 650898 57206 651134
rect 87690 651218 87926 651454
rect 87690 650898 87926 651134
rect 118410 651218 118646 651454
rect 118410 650898 118646 651134
rect 149130 651218 149366 651454
rect 149130 650898 149366 651134
rect 179850 651218 180086 651454
rect 179850 650898 180086 651134
rect 210570 651218 210806 651454
rect 210570 650898 210806 651134
rect 241290 651218 241526 651454
rect 241290 650898 241526 651134
rect 272010 651218 272246 651454
rect 272010 650898 272246 651134
rect 302730 651218 302966 651454
rect 302730 650898 302966 651134
rect 333450 651218 333686 651454
rect 333450 650898 333686 651134
rect 364170 651218 364406 651454
rect 364170 650898 364406 651134
rect 394890 651218 395126 651454
rect 394890 650898 395126 651134
rect 425610 651218 425846 651454
rect 425610 650898 425846 651134
rect 456330 651218 456566 651454
rect 456330 650898 456566 651134
rect 487050 651218 487286 651454
rect 487050 650898 487286 651134
rect 517770 651218 518006 651454
rect 517770 650898 518006 651134
rect 548490 651218 548726 651454
rect 548490 650898 548726 651134
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 41610 618938 41846 619174
rect 41610 618618 41846 618854
rect 72330 618938 72566 619174
rect 72330 618618 72566 618854
rect 103050 618938 103286 619174
rect 103050 618618 103286 618854
rect 133770 618938 134006 619174
rect 133770 618618 134006 618854
rect 164490 618938 164726 619174
rect 164490 618618 164726 618854
rect 195210 618938 195446 619174
rect 195210 618618 195446 618854
rect 225930 618938 226166 619174
rect 225930 618618 226166 618854
rect 256650 618938 256886 619174
rect 256650 618618 256886 618854
rect 287370 618938 287606 619174
rect 287370 618618 287606 618854
rect 318090 618938 318326 619174
rect 318090 618618 318326 618854
rect 348810 618938 349046 619174
rect 348810 618618 349046 618854
rect 379530 618938 379766 619174
rect 379530 618618 379766 618854
rect 410250 618938 410486 619174
rect 410250 618618 410486 618854
rect 440970 618938 441206 619174
rect 440970 618618 441206 618854
rect 471690 618938 471926 619174
rect 471690 618618 471926 618854
rect 502410 618938 502646 619174
rect 502410 618618 502646 618854
rect 533130 618938 533366 619174
rect 533130 618618 533366 618854
rect 26250 615218 26486 615454
rect 26250 614898 26486 615134
rect 56970 615218 57206 615454
rect 56970 614898 57206 615134
rect 87690 615218 87926 615454
rect 87690 614898 87926 615134
rect 118410 615218 118646 615454
rect 118410 614898 118646 615134
rect 149130 615218 149366 615454
rect 149130 614898 149366 615134
rect 179850 615218 180086 615454
rect 179850 614898 180086 615134
rect 210570 615218 210806 615454
rect 210570 614898 210806 615134
rect 241290 615218 241526 615454
rect 241290 614898 241526 615134
rect 272010 615218 272246 615454
rect 272010 614898 272246 615134
rect 302730 615218 302966 615454
rect 302730 614898 302966 615134
rect 333450 615218 333686 615454
rect 333450 614898 333686 615134
rect 364170 615218 364406 615454
rect 364170 614898 364406 615134
rect 394890 615218 395126 615454
rect 394890 614898 395126 615134
rect 425610 615218 425846 615454
rect 425610 614898 425846 615134
rect 456330 615218 456566 615454
rect 456330 614898 456566 615134
rect 487050 615218 487286 615454
rect 487050 614898 487286 615134
rect 517770 615218 518006 615454
rect 517770 614898 518006 615134
rect 548490 615218 548726 615454
rect 548490 614898 548726 615134
rect 24146 601538 24382 601774
rect 24466 601538 24702 601774
rect 24146 601218 24382 601454
rect 24466 601218 24702 601454
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 41610 582938 41846 583174
rect 41610 582618 41846 582854
rect 72330 582938 72566 583174
rect 72330 582618 72566 582854
rect 103050 582938 103286 583174
rect 103050 582618 103286 582854
rect 133770 582938 134006 583174
rect 133770 582618 134006 582854
rect 164490 582938 164726 583174
rect 164490 582618 164726 582854
rect 195210 582938 195446 583174
rect 195210 582618 195446 582854
rect 225930 582938 226166 583174
rect 225930 582618 226166 582854
rect 256650 582938 256886 583174
rect 256650 582618 256886 582854
rect 287370 582938 287606 583174
rect 287370 582618 287606 582854
rect 318090 582938 318326 583174
rect 318090 582618 318326 582854
rect 348810 582938 349046 583174
rect 348810 582618 349046 582854
rect 379530 582938 379766 583174
rect 379530 582618 379766 582854
rect 410250 582938 410486 583174
rect 410250 582618 410486 582854
rect 440970 582938 441206 583174
rect 440970 582618 441206 582854
rect 471690 582938 471926 583174
rect 471690 582618 471926 582854
rect 502410 582938 502646 583174
rect 502410 582618 502646 582854
rect 533130 582938 533366 583174
rect 533130 582618 533366 582854
rect 26250 579218 26486 579454
rect 26250 578898 26486 579134
rect 56970 579218 57206 579454
rect 56970 578898 57206 579134
rect 87690 579218 87926 579454
rect 87690 578898 87926 579134
rect 118410 579218 118646 579454
rect 118410 578898 118646 579134
rect 149130 579218 149366 579454
rect 149130 578898 149366 579134
rect 179850 579218 180086 579454
rect 179850 578898 180086 579134
rect 210570 579218 210806 579454
rect 210570 578898 210806 579134
rect 241290 579218 241526 579454
rect 241290 578898 241526 579134
rect 272010 579218 272246 579454
rect 272010 578898 272246 579134
rect 302730 579218 302966 579454
rect 302730 578898 302966 579134
rect 333450 579218 333686 579454
rect 333450 578898 333686 579134
rect 364170 579218 364406 579454
rect 364170 578898 364406 579134
rect 394890 579218 395126 579454
rect 394890 578898 395126 579134
rect 425610 579218 425846 579454
rect 425610 578898 425846 579134
rect 456330 579218 456566 579454
rect 456330 578898 456566 579134
rect 487050 579218 487286 579454
rect 487050 578898 487286 579134
rect 517770 579218 518006 579454
rect 517770 578898 518006 579134
rect 548490 579218 548726 579454
rect 548490 578898 548726 579134
rect 24146 565538 24382 565774
rect 24466 565538 24702 565774
rect 24146 565218 24382 565454
rect 24466 565218 24702 565454
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 41610 546938 41846 547174
rect 41610 546618 41846 546854
rect 72330 546938 72566 547174
rect 72330 546618 72566 546854
rect 103050 546938 103286 547174
rect 103050 546618 103286 546854
rect 133770 546938 134006 547174
rect 133770 546618 134006 546854
rect 164490 546938 164726 547174
rect 164490 546618 164726 546854
rect 195210 546938 195446 547174
rect 195210 546618 195446 546854
rect 225930 546938 226166 547174
rect 225930 546618 226166 546854
rect 256650 546938 256886 547174
rect 256650 546618 256886 546854
rect 287370 546938 287606 547174
rect 287370 546618 287606 546854
rect 318090 546938 318326 547174
rect 318090 546618 318326 546854
rect 348810 546938 349046 547174
rect 348810 546618 349046 546854
rect 379530 546938 379766 547174
rect 379530 546618 379766 546854
rect 410250 546938 410486 547174
rect 410250 546618 410486 546854
rect 440970 546938 441206 547174
rect 440970 546618 441206 546854
rect 471690 546938 471926 547174
rect 471690 546618 471926 546854
rect 502410 546938 502646 547174
rect 502410 546618 502646 546854
rect 533130 546938 533366 547174
rect 533130 546618 533366 546854
rect 26250 543218 26486 543454
rect 26250 542898 26486 543134
rect 56970 543218 57206 543454
rect 56970 542898 57206 543134
rect 87690 543218 87926 543454
rect 87690 542898 87926 543134
rect 118410 543218 118646 543454
rect 118410 542898 118646 543134
rect 149130 543218 149366 543454
rect 149130 542898 149366 543134
rect 179850 543218 180086 543454
rect 179850 542898 180086 543134
rect 210570 543218 210806 543454
rect 210570 542898 210806 543134
rect 241290 543218 241526 543454
rect 241290 542898 241526 543134
rect 272010 543218 272246 543454
rect 272010 542898 272246 543134
rect 302730 543218 302966 543454
rect 302730 542898 302966 543134
rect 333450 543218 333686 543454
rect 333450 542898 333686 543134
rect 364170 543218 364406 543454
rect 364170 542898 364406 543134
rect 394890 543218 395126 543454
rect 394890 542898 395126 543134
rect 425610 543218 425846 543454
rect 425610 542898 425846 543134
rect 456330 543218 456566 543454
rect 456330 542898 456566 543134
rect 487050 543218 487286 543454
rect 487050 542898 487286 543134
rect 517770 543218 518006 543454
rect 517770 542898 518006 543134
rect 548490 543218 548726 543454
rect 548490 542898 548726 543134
rect 24146 529538 24382 529774
rect 24466 529538 24702 529774
rect 24146 529218 24382 529454
rect 24466 529218 24702 529454
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 41610 510938 41846 511174
rect 41610 510618 41846 510854
rect 72330 510938 72566 511174
rect 72330 510618 72566 510854
rect 103050 510938 103286 511174
rect 103050 510618 103286 510854
rect 133770 510938 134006 511174
rect 133770 510618 134006 510854
rect 164490 510938 164726 511174
rect 164490 510618 164726 510854
rect 195210 510938 195446 511174
rect 195210 510618 195446 510854
rect 225930 510938 226166 511174
rect 225930 510618 226166 510854
rect 256650 510938 256886 511174
rect 256650 510618 256886 510854
rect 287370 510938 287606 511174
rect 287370 510618 287606 510854
rect 318090 510938 318326 511174
rect 318090 510618 318326 510854
rect 348810 510938 349046 511174
rect 348810 510618 349046 510854
rect 379530 510938 379766 511174
rect 379530 510618 379766 510854
rect 410250 510938 410486 511174
rect 410250 510618 410486 510854
rect 440970 510938 441206 511174
rect 440970 510618 441206 510854
rect 471690 510938 471926 511174
rect 471690 510618 471926 510854
rect 502410 510938 502646 511174
rect 502410 510618 502646 510854
rect 533130 510938 533366 511174
rect 533130 510618 533366 510854
rect 26250 507218 26486 507454
rect 26250 506898 26486 507134
rect 56970 507218 57206 507454
rect 56970 506898 57206 507134
rect 87690 507218 87926 507454
rect 87690 506898 87926 507134
rect 118410 507218 118646 507454
rect 118410 506898 118646 507134
rect 149130 507218 149366 507454
rect 149130 506898 149366 507134
rect 179850 507218 180086 507454
rect 179850 506898 180086 507134
rect 210570 507218 210806 507454
rect 210570 506898 210806 507134
rect 241290 507218 241526 507454
rect 241290 506898 241526 507134
rect 272010 507218 272246 507454
rect 272010 506898 272246 507134
rect 302730 507218 302966 507454
rect 302730 506898 302966 507134
rect 333450 507218 333686 507454
rect 333450 506898 333686 507134
rect 364170 507218 364406 507454
rect 364170 506898 364406 507134
rect 394890 507218 395126 507454
rect 394890 506898 395126 507134
rect 425610 507218 425846 507454
rect 425610 506898 425846 507134
rect 456330 507218 456566 507454
rect 456330 506898 456566 507134
rect 487050 507218 487286 507454
rect 487050 506898 487286 507134
rect 517770 507218 518006 507454
rect 517770 506898 518006 507134
rect 548490 507218 548726 507454
rect 548490 506898 548726 507134
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 41610 474938 41846 475174
rect 41610 474618 41846 474854
rect 72330 474938 72566 475174
rect 72330 474618 72566 474854
rect 103050 474938 103286 475174
rect 103050 474618 103286 474854
rect 133770 474938 134006 475174
rect 133770 474618 134006 474854
rect 164490 474938 164726 475174
rect 164490 474618 164726 474854
rect 195210 474938 195446 475174
rect 195210 474618 195446 474854
rect 225930 474938 226166 475174
rect 225930 474618 226166 474854
rect 256650 474938 256886 475174
rect 256650 474618 256886 474854
rect 287370 474938 287606 475174
rect 287370 474618 287606 474854
rect 318090 474938 318326 475174
rect 318090 474618 318326 474854
rect 348810 474938 349046 475174
rect 348810 474618 349046 474854
rect 379530 474938 379766 475174
rect 379530 474618 379766 474854
rect 410250 474938 410486 475174
rect 410250 474618 410486 474854
rect 440970 474938 441206 475174
rect 440970 474618 441206 474854
rect 471690 474938 471926 475174
rect 471690 474618 471926 474854
rect 502410 474938 502646 475174
rect 502410 474618 502646 474854
rect 533130 474938 533366 475174
rect 533130 474618 533366 474854
rect 26250 471218 26486 471454
rect 26250 470898 26486 471134
rect 56970 471218 57206 471454
rect 56970 470898 57206 471134
rect 87690 471218 87926 471454
rect 87690 470898 87926 471134
rect 118410 471218 118646 471454
rect 118410 470898 118646 471134
rect 149130 471218 149366 471454
rect 149130 470898 149366 471134
rect 179850 471218 180086 471454
rect 179850 470898 180086 471134
rect 210570 471218 210806 471454
rect 210570 470898 210806 471134
rect 241290 471218 241526 471454
rect 241290 470898 241526 471134
rect 272010 471218 272246 471454
rect 272010 470898 272246 471134
rect 302730 471218 302966 471454
rect 302730 470898 302966 471134
rect 333450 471218 333686 471454
rect 333450 470898 333686 471134
rect 364170 471218 364406 471454
rect 364170 470898 364406 471134
rect 394890 471218 395126 471454
rect 394890 470898 395126 471134
rect 425610 471218 425846 471454
rect 425610 470898 425846 471134
rect 456330 471218 456566 471454
rect 456330 470898 456566 471134
rect 487050 471218 487286 471454
rect 487050 470898 487286 471134
rect 517770 471218 518006 471454
rect 517770 470898 518006 471134
rect 548490 471218 548726 471454
rect 548490 470898 548726 471134
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 41610 438938 41846 439174
rect 41610 438618 41846 438854
rect 72330 438938 72566 439174
rect 72330 438618 72566 438854
rect 103050 438938 103286 439174
rect 103050 438618 103286 438854
rect 133770 438938 134006 439174
rect 133770 438618 134006 438854
rect 164490 438938 164726 439174
rect 164490 438618 164726 438854
rect 195210 438938 195446 439174
rect 195210 438618 195446 438854
rect 225930 438938 226166 439174
rect 225930 438618 226166 438854
rect 256650 438938 256886 439174
rect 256650 438618 256886 438854
rect 287370 438938 287606 439174
rect 287370 438618 287606 438854
rect 318090 438938 318326 439174
rect 318090 438618 318326 438854
rect 348810 438938 349046 439174
rect 348810 438618 349046 438854
rect 379530 438938 379766 439174
rect 379530 438618 379766 438854
rect 410250 438938 410486 439174
rect 410250 438618 410486 438854
rect 440970 438938 441206 439174
rect 440970 438618 441206 438854
rect 471690 438938 471926 439174
rect 471690 438618 471926 438854
rect 502410 438938 502646 439174
rect 502410 438618 502646 438854
rect 533130 438938 533366 439174
rect 533130 438618 533366 438854
rect 26250 435218 26486 435454
rect 26250 434898 26486 435134
rect 56970 435218 57206 435454
rect 56970 434898 57206 435134
rect 87690 435218 87926 435454
rect 87690 434898 87926 435134
rect 118410 435218 118646 435454
rect 118410 434898 118646 435134
rect 149130 435218 149366 435454
rect 149130 434898 149366 435134
rect 179850 435218 180086 435454
rect 179850 434898 180086 435134
rect 210570 435218 210806 435454
rect 210570 434898 210806 435134
rect 241290 435218 241526 435454
rect 241290 434898 241526 435134
rect 272010 435218 272246 435454
rect 272010 434898 272246 435134
rect 302730 435218 302966 435454
rect 302730 434898 302966 435134
rect 333450 435218 333686 435454
rect 333450 434898 333686 435134
rect 364170 435218 364406 435454
rect 364170 434898 364406 435134
rect 394890 435218 395126 435454
rect 394890 434898 395126 435134
rect 425610 435218 425846 435454
rect 425610 434898 425846 435134
rect 456330 435218 456566 435454
rect 456330 434898 456566 435134
rect 487050 435218 487286 435454
rect 487050 434898 487286 435134
rect 517770 435218 518006 435454
rect 517770 434898 518006 435134
rect 548490 435218 548726 435454
rect 548490 434898 548726 435134
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 41610 402938 41846 403174
rect 41610 402618 41846 402854
rect 72330 402938 72566 403174
rect 72330 402618 72566 402854
rect 103050 402938 103286 403174
rect 103050 402618 103286 402854
rect 133770 402938 134006 403174
rect 133770 402618 134006 402854
rect 164490 402938 164726 403174
rect 164490 402618 164726 402854
rect 195210 402938 195446 403174
rect 195210 402618 195446 402854
rect 225930 402938 226166 403174
rect 225930 402618 226166 402854
rect 256650 402938 256886 403174
rect 256650 402618 256886 402854
rect 287370 402938 287606 403174
rect 287370 402618 287606 402854
rect 318090 402938 318326 403174
rect 318090 402618 318326 402854
rect 348810 402938 349046 403174
rect 348810 402618 349046 402854
rect 379530 402938 379766 403174
rect 379530 402618 379766 402854
rect 410250 402938 410486 403174
rect 410250 402618 410486 402854
rect 440970 402938 441206 403174
rect 440970 402618 441206 402854
rect 471690 402938 471926 403174
rect 471690 402618 471926 402854
rect 502410 402938 502646 403174
rect 502410 402618 502646 402854
rect 533130 402938 533366 403174
rect 533130 402618 533366 402854
rect 26250 399218 26486 399454
rect 26250 398898 26486 399134
rect 56970 399218 57206 399454
rect 56970 398898 57206 399134
rect 87690 399218 87926 399454
rect 87690 398898 87926 399134
rect 118410 399218 118646 399454
rect 118410 398898 118646 399134
rect 149130 399218 149366 399454
rect 149130 398898 149366 399134
rect 179850 399218 180086 399454
rect 179850 398898 180086 399134
rect 210570 399218 210806 399454
rect 210570 398898 210806 399134
rect 241290 399218 241526 399454
rect 241290 398898 241526 399134
rect 272010 399218 272246 399454
rect 272010 398898 272246 399134
rect 302730 399218 302966 399454
rect 302730 398898 302966 399134
rect 333450 399218 333686 399454
rect 333450 398898 333686 399134
rect 364170 399218 364406 399454
rect 364170 398898 364406 399134
rect 394890 399218 395126 399454
rect 394890 398898 395126 399134
rect 425610 399218 425846 399454
rect 425610 398898 425846 399134
rect 456330 399218 456566 399454
rect 456330 398898 456566 399134
rect 487050 399218 487286 399454
rect 487050 398898 487286 399134
rect 517770 399218 518006 399454
rect 517770 398898 518006 399134
rect 548490 399218 548726 399454
rect 548490 398898 548726 399134
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 41610 366938 41846 367174
rect 41610 366618 41846 366854
rect 72330 366938 72566 367174
rect 72330 366618 72566 366854
rect 103050 366938 103286 367174
rect 103050 366618 103286 366854
rect 133770 366938 134006 367174
rect 133770 366618 134006 366854
rect 164490 366938 164726 367174
rect 164490 366618 164726 366854
rect 195210 366938 195446 367174
rect 195210 366618 195446 366854
rect 225930 366938 226166 367174
rect 225930 366618 226166 366854
rect 256650 366938 256886 367174
rect 256650 366618 256886 366854
rect 287370 366938 287606 367174
rect 287370 366618 287606 366854
rect 318090 366938 318326 367174
rect 318090 366618 318326 366854
rect 348810 366938 349046 367174
rect 348810 366618 349046 366854
rect 379530 366938 379766 367174
rect 379530 366618 379766 366854
rect 410250 366938 410486 367174
rect 410250 366618 410486 366854
rect 440970 366938 441206 367174
rect 440970 366618 441206 366854
rect 471690 366938 471926 367174
rect 471690 366618 471926 366854
rect 502410 366938 502646 367174
rect 502410 366618 502646 366854
rect 533130 366938 533366 367174
rect 533130 366618 533366 366854
rect 26250 363218 26486 363454
rect 26250 362898 26486 363134
rect 56970 363218 57206 363454
rect 56970 362898 57206 363134
rect 87690 363218 87926 363454
rect 87690 362898 87926 363134
rect 118410 363218 118646 363454
rect 118410 362898 118646 363134
rect 149130 363218 149366 363454
rect 149130 362898 149366 363134
rect 179850 363218 180086 363454
rect 179850 362898 180086 363134
rect 210570 363218 210806 363454
rect 210570 362898 210806 363134
rect 241290 363218 241526 363454
rect 241290 362898 241526 363134
rect 272010 363218 272246 363454
rect 272010 362898 272246 363134
rect 302730 363218 302966 363454
rect 302730 362898 302966 363134
rect 333450 363218 333686 363454
rect 333450 362898 333686 363134
rect 364170 363218 364406 363454
rect 364170 362898 364406 363134
rect 394890 363218 395126 363454
rect 394890 362898 395126 363134
rect 425610 363218 425846 363454
rect 425610 362898 425846 363134
rect 456330 363218 456566 363454
rect 456330 362898 456566 363134
rect 487050 363218 487286 363454
rect 487050 362898 487286 363134
rect 517770 363218 518006 363454
rect 517770 362898 518006 363134
rect 548490 363218 548726 363454
rect 548490 362898 548726 363134
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 41610 330938 41846 331174
rect 41610 330618 41846 330854
rect 72330 330938 72566 331174
rect 72330 330618 72566 330854
rect 103050 330938 103286 331174
rect 103050 330618 103286 330854
rect 133770 330938 134006 331174
rect 133770 330618 134006 330854
rect 164490 330938 164726 331174
rect 164490 330618 164726 330854
rect 195210 330938 195446 331174
rect 195210 330618 195446 330854
rect 225930 330938 226166 331174
rect 225930 330618 226166 330854
rect 256650 330938 256886 331174
rect 256650 330618 256886 330854
rect 287370 330938 287606 331174
rect 287370 330618 287606 330854
rect 318090 330938 318326 331174
rect 318090 330618 318326 330854
rect 348810 330938 349046 331174
rect 348810 330618 349046 330854
rect 379530 330938 379766 331174
rect 379530 330618 379766 330854
rect 410250 330938 410486 331174
rect 410250 330618 410486 330854
rect 440970 330938 441206 331174
rect 440970 330618 441206 330854
rect 471690 330938 471926 331174
rect 471690 330618 471926 330854
rect 502410 330938 502646 331174
rect 502410 330618 502646 330854
rect 533130 330938 533366 331174
rect 533130 330618 533366 330854
rect 26250 327218 26486 327454
rect 26250 326898 26486 327134
rect 56970 327218 57206 327454
rect 56970 326898 57206 327134
rect 87690 327218 87926 327454
rect 87690 326898 87926 327134
rect 118410 327218 118646 327454
rect 118410 326898 118646 327134
rect 149130 327218 149366 327454
rect 149130 326898 149366 327134
rect 179850 327218 180086 327454
rect 179850 326898 180086 327134
rect 210570 327218 210806 327454
rect 210570 326898 210806 327134
rect 241290 327218 241526 327454
rect 241290 326898 241526 327134
rect 272010 327218 272246 327454
rect 272010 326898 272246 327134
rect 302730 327218 302966 327454
rect 302730 326898 302966 327134
rect 333450 327218 333686 327454
rect 333450 326898 333686 327134
rect 364170 327218 364406 327454
rect 364170 326898 364406 327134
rect 394890 327218 395126 327454
rect 394890 326898 395126 327134
rect 425610 327218 425846 327454
rect 425610 326898 425846 327134
rect 456330 327218 456566 327454
rect 456330 326898 456566 327134
rect 487050 327218 487286 327454
rect 487050 326898 487286 327134
rect 517770 327218 518006 327454
rect 517770 326898 518006 327134
rect 548490 327218 548726 327454
rect 548490 326898 548726 327134
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 41610 294938 41846 295174
rect 41610 294618 41846 294854
rect 72330 294938 72566 295174
rect 72330 294618 72566 294854
rect 103050 294938 103286 295174
rect 103050 294618 103286 294854
rect 133770 294938 134006 295174
rect 133770 294618 134006 294854
rect 164490 294938 164726 295174
rect 164490 294618 164726 294854
rect 195210 294938 195446 295174
rect 195210 294618 195446 294854
rect 225930 294938 226166 295174
rect 225930 294618 226166 294854
rect 256650 294938 256886 295174
rect 256650 294618 256886 294854
rect 287370 294938 287606 295174
rect 287370 294618 287606 294854
rect 318090 294938 318326 295174
rect 318090 294618 318326 294854
rect 348810 294938 349046 295174
rect 348810 294618 349046 294854
rect 379530 294938 379766 295174
rect 379530 294618 379766 294854
rect 410250 294938 410486 295174
rect 410250 294618 410486 294854
rect 440970 294938 441206 295174
rect 440970 294618 441206 294854
rect 471690 294938 471926 295174
rect 471690 294618 471926 294854
rect 502410 294938 502646 295174
rect 502410 294618 502646 294854
rect 533130 294938 533366 295174
rect 533130 294618 533366 294854
rect 26250 291218 26486 291454
rect 26250 290898 26486 291134
rect 56970 291218 57206 291454
rect 56970 290898 57206 291134
rect 87690 291218 87926 291454
rect 87690 290898 87926 291134
rect 118410 291218 118646 291454
rect 118410 290898 118646 291134
rect 149130 291218 149366 291454
rect 149130 290898 149366 291134
rect 179850 291218 180086 291454
rect 179850 290898 180086 291134
rect 210570 291218 210806 291454
rect 210570 290898 210806 291134
rect 241290 291218 241526 291454
rect 241290 290898 241526 291134
rect 272010 291218 272246 291454
rect 272010 290898 272246 291134
rect 302730 291218 302966 291454
rect 302730 290898 302966 291134
rect 333450 291218 333686 291454
rect 333450 290898 333686 291134
rect 364170 291218 364406 291454
rect 364170 290898 364406 291134
rect 394890 291218 395126 291454
rect 394890 290898 395126 291134
rect 425610 291218 425846 291454
rect 425610 290898 425846 291134
rect 456330 291218 456566 291454
rect 456330 290898 456566 291134
rect 487050 291218 487286 291454
rect 487050 290898 487286 291134
rect 517770 291218 518006 291454
rect 517770 290898 518006 291134
rect 548490 291218 548726 291454
rect 548490 290898 548726 291134
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 41610 258938 41846 259174
rect 41610 258618 41846 258854
rect 72330 258938 72566 259174
rect 72330 258618 72566 258854
rect 103050 258938 103286 259174
rect 103050 258618 103286 258854
rect 133770 258938 134006 259174
rect 133770 258618 134006 258854
rect 164490 258938 164726 259174
rect 164490 258618 164726 258854
rect 195210 258938 195446 259174
rect 195210 258618 195446 258854
rect 225930 258938 226166 259174
rect 225930 258618 226166 258854
rect 256650 258938 256886 259174
rect 256650 258618 256886 258854
rect 287370 258938 287606 259174
rect 287370 258618 287606 258854
rect 318090 258938 318326 259174
rect 318090 258618 318326 258854
rect 348810 258938 349046 259174
rect 348810 258618 349046 258854
rect 379530 258938 379766 259174
rect 379530 258618 379766 258854
rect 410250 258938 410486 259174
rect 410250 258618 410486 258854
rect 440970 258938 441206 259174
rect 440970 258618 441206 258854
rect 471690 258938 471926 259174
rect 471690 258618 471926 258854
rect 502410 258938 502646 259174
rect 502410 258618 502646 258854
rect 533130 258938 533366 259174
rect 533130 258618 533366 258854
rect 26250 255218 26486 255454
rect 26250 254898 26486 255134
rect 56970 255218 57206 255454
rect 56970 254898 57206 255134
rect 87690 255218 87926 255454
rect 87690 254898 87926 255134
rect 118410 255218 118646 255454
rect 118410 254898 118646 255134
rect 149130 255218 149366 255454
rect 149130 254898 149366 255134
rect 179850 255218 180086 255454
rect 179850 254898 180086 255134
rect 210570 255218 210806 255454
rect 210570 254898 210806 255134
rect 241290 255218 241526 255454
rect 241290 254898 241526 255134
rect 272010 255218 272246 255454
rect 272010 254898 272246 255134
rect 302730 255218 302966 255454
rect 302730 254898 302966 255134
rect 333450 255218 333686 255454
rect 333450 254898 333686 255134
rect 364170 255218 364406 255454
rect 364170 254898 364406 255134
rect 394890 255218 395126 255454
rect 394890 254898 395126 255134
rect 425610 255218 425846 255454
rect 425610 254898 425846 255134
rect 456330 255218 456566 255454
rect 456330 254898 456566 255134
rect 487050 255218 487286 255454
rect 487050 254898 487286 255134
rect 517770 255218 518006 255454
rect 517770 254898 518006 255134
rect 548490 255218 548726 255454
rect 548490 254898 548726 255134
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 41610 222938 41846 223174
rect 41610 222618 41846 222854
rect 72330 222938 72566 223174
rect 72330 222618 72566 222854
rect 103050 222938 103286 223174
rect 103050 222618 103286 222854
rect 133770 222938 134006 223174
rect 133770 222618 134006 222854
rect 164490 222938 164726 223174
rect 164490 222618 164726 222854
rect 195210 222938 195446 223174
rect 195210 222618 195446 222854
rect 225930 222938 226166 223174
rect 225930 222618 226166 222854
rect 256650 222938 256886 223174
rect 256650 222618 256886 222854
rect 287370 222938 287606 223174
rect 287370 222618 287606 222854
rect 318090 222938 318326 223174
rect 318090 222618 318326 222854
rect 348810 222938 349046 223174
rect 348810 222618 349046 222854
rect 379530 222938 379766 223174
rect 379530 222618 379766 222854
rect 410250 222938 410486 223174
rect 410250 222618 410486 222854
rect 440970 222938 441206 223174
rect 440970 222618 441206 222854
rect 471690 222938 471926 223174
rect 471690 222618 471926 222854
rect 502410 222938 502646 223174
rect 502410 222618 502646 222854
rect 533130 222938 533366 223174
rect 533130 222618 533366 222854
rect 26250 219218 26486 219454
rect 26250 218898 26486 219134
rect 56970 219218 57206 219454
rect 56970 218898 57206 219134
rect 87690 219218 87926 219454
rect 87690 218898 87926 219134
rect 118410 219218 118646 219454
rect 118410 218898 118646 219134
rect 149130 219218 149366 219454
rect 149130 218898 149366 219134
rect 179850 219218 180086 219454
rect 179850 218898 180086 219134
rect 210570 219218 210806 219454
rect 210570 218898 210806 219134
rect 241290 219218 241526 219454
rect 241290 218898 241526 219134
rect 272010 219218 272246 219454
rect 272010 218898 272246 219134
rect 302730 219218 302966 219454
rect 302730 218898 302966 219134
rect 333450 219218 333686 219454
rect 333450 218898 333686 219134
rect 364170 219218 364406 219454
rect 364170 218898 364406 219134
rect 394890 219218 395126 219454
rect 394890 218898 395126 219134
rect 425610 219218 425846 219454
rect 425610 218898 425846 219134
rect 456330 219218 456566 219454
rect 456330 218898 456566 219134
rect 487050 219218 487286 219454
rect 487050 218898 487286 219134
rect 517770 219218 518006 219454
rect 517770 218898 518006 219134
rect 548490 219218 548726 219454
rect 548490 218898 548726 219134
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 41610 186938 41846 187174
rect 41610 186618 41846 186854
rect 72330 186938 72566 187174
rect 72330 186618 72566 186854
rect 103050 186938 103286 187174
rect 103050 186618 103286 186854
rect 133770 186938 134006 187174
rect 133770 186618 134006 186854
rect 164490 186938 164726 187174
rect 164490 186618 164726 186854
rect 195210 186938 195446 187174
rect 195210 186618 195446 186854
rect 225930 186938 226166 187174
rect 225930 186618 226166 186854
rect 256650 186938 256886 187174
rect 256650 186618 256886 186854
rect 287370 186938 287606 187174
rect 287370 186618 287606 186854
rect 318090 186938 318326 187174
rect 318090 186618 318326 186854
rect 348810 186938 349046 187174
rect 348810 186618 349046 186854
rect 379530 186938 379766 187174
rect 379530 186618 379766 186854
rect 410250 186938 410486 187174
rect 410250 186618 410486 186854
rect 440970 186938 441206 187174
rect 440970 186618 441206 186854
rect 471690 186938 471926 187174
rect 471690 186618 471926 186854
rect 502410 186938 502646 187174
rect 502410 186618 502646 186854
rect 533130 186938 533366 187174
rect 533130 186618 533366 186854
rect 26250 183218 26486 183454
rect 26250 182898 26486 183134
rect 56970 183218 57206 183454
rect 56970 182898 57206 183134
rect 87690 183218 87926 183454
rect 87690 182898 87926 183134
rect 118410 183218 118646 183454
rect 118410 182898 118646 183134
rect 149130 183218 149366 183454
rect 149130 182898 149366 183134
rect 179850 183218 180086 183454
rect 179850 182898 180086 183134
rect 210570 183218 210806 183454
rect 210570 182898 210806 183134
rect 241290 183218 241526 183454
rect 241290 182898 241526 183134
rect 272010 183218 272246 183454
rect 272010 182898 272246 183134
rect 302730 183218 302966 183454
rect 302730 182898 302966 183134
rect 333450 183218 333686 183454
rect 333450 182898 333686 183134
rect 364170 183218 364406 183454
rect 364170 182898 364406 183134
rect 394890 183218 395126 183454
rect 394890 182898 395126 183134
rect 425610 183218 425846 183454
rect 425610 182898 425846 183134
rect 456330 183218 456566 183454
rect 456330 182898 456566 183134
rect 487050 183218 487286 183454
rect 487050 182898 487286 183134
rect 517770 183218 518006 183454
rect 517770 182898 518006 183134
rect 548490 183218 548726 183454
rect 548490 182898 548726 183134
rect 24146 169538 24382 169774
rect 24466 169538 24702 169774
rect 24146 169218 24382 169454
rect 24466 169218 24702 169454
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 41610 150938 41846 151174
rect 41610 150618 41846 150854
rect 72330 150938 72566 151174
rect 72330 150618 72566 150854
rect 103050 150938 103286 151174
rect 103050 150618 103286 150854
rect 133770 150938 134006 151174
rect 133770 150618 134006 150854
rect 164490 150938 164726 151174
rect 164490 150618 164726 150854
rect 195210 150938 195446 151174
rect 195210 150618 195446 150854
rect 225930 150938 226166 151174
rect 225930 150618 226166 150854
rect 256650 150938 256886 151174
rect 256650 150618 256886 150854
rect 287370 150938 287606 151174
rect 287370 150618 287606 150854
rect 318090 150938 318326 151174
rect 318090 150618 318326 150854
rect 348810 150938 349046 151174
rect 348810 150618 349046 150854
rect 379530 150938 379766 151174
rect 379530 150618 379766 150854
rect 410250 150938 410486 151174
rect 410250 150618 410486 150854
rect 440970 150938 441206 151174
rect 440970 150618 441206 150854
rect 471690 150938 471926 151174
rect 471690 150618 471926 150854
rect 502410 150938 502646 151174
rect 502410 150618 502646 150854
rect 533130 150938 533366 151174
rect 533130 150618 533366 150854
rect 26250 147218 26486 147454
rect 26250 146898 26486 147134
rect 56970 147218 57206 147454
rect 56970 146898 57206 147134
rect 87690 147218 87926 147454
rect 87690 146898 87926 147134
rect 118410 147218 118646 147454
rect 118410 146898 118646 147134
rect 149130 147218 149366 147454
rect 149130 146898 149366 147134
rect 179850 147218 180086 147454
rect 179850 146898 180086 147134
rect 210570 147218 210806 147454
rect 210570 146898 210806 147134
rect 241290 147218 241526 147454
rect 241290 146898 241526 147134
rect 272010 147218 272246 147454
rect 272010 146898 272246 147134
rect 302730 147218 302966 147454
rect 302730 146898 302966 147134
rect 333450 147218 333686 147454
rect 333450 146898 333686 147134
rect 364170 147218 364406 147454
rect 364170 146898 364406 147134
rect 394890 147218 395126 147454
rect 394890 146898 395126 147134
rect 425610 147218 425846 147454
rect 425610 146898 425846 147134
rect 456330 147218 456566 147454
rect 456330 146898 456566 147134
rect 487050 147218 487286 147454
rect 487050 146898 487286 147134
rect 517770 147218 518006 147454
rect 517770 146898 518006 147134
rect 548490 147218 548726 147454
rect 548490 146898 548726 147134
rect 24146 133538 24382 133774
rect 24466 133538 24702 133774
rect 24146 133218 24382 133454
rect 24466 133218 24702 133454
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 41610 114938 41846 115174
rect 41610 114618 41846 114854
rect 72330 114938 72566 115174
rect 72330 114618 72566 114854
rect 103050 114938 103286 115174
rect 103050 114618 103286 114854
rect 133770 114938 134006 115174
rect 133770 114618 134006 114854
rect 164490 114938 164726 115174
rect 164490 114618 164726 114854
rect 195210 114938 195446 115174
rect 195210 114618 195446 114854
rect 225930 114938 226166 115174
rect 225930 114618 226166 114854
rect 256650 114938 256886 115174
rect 256650 114618 256886 114854
rect 287370 114938 287606 115174
rect 287370 114618 287606 114854
rect 318090 114938 318326 115174
rect 318090 114618 318326 114854
rect 348810 114938 349046 115174
rect 348810 114618 349046 114854
rect 379530 114938 379766 115174
rect 379530 114618 379766 114854
rect 410250 114938 410486 115174
rect 410250 114618 410486 114854
rect 440970 114938 441206 115174
rect 440970 114618 441206 114854
rect 471690 114938 471926 115174
rect 471690 114618 471926 114854
rect 502410 114938 502646 115174
rect 502410 114618 502646 114854
rect 533130 114938 533366 115174
rect 533130 114618 533366 114854
rect 26250 111218 26486 111454
rect 26250 110898 26486 111134
rect 56970 111218 57206 111454
rect 56970 110898 57206 111134
rect 87690 111218 87926 111454
rect 87690 110898 87926 111134
rect 118410 111218 118646 111454
rect 118410 110898 118646 111134
rect 149130 111218 149366 111454
rect 149130 110898 149366 111134
rect 179850 111218 180086 111454
rect 179850 110898 180086 111134
rect 210570 111218 210806 111454
rect 210570 110898 210806 111134
rect 241290 111218 241526 111454
rect 241290 110898 241526 111134
rect 272010 111218 272246 111454
rect 272010 110898 272246 111134
rect 302730 111218 302966 111454
rect 302730 110898 302966 111134
rect 333450 111218 333686 111454
rect 333450 110898 333686 111134
rect 364170 111218 364406 111454
rect 364170 110898 364406 111134
rect 394890 111218 395126 111454
rect 394890 110898 395126 111134
rect 425610 111218 425846 111454
rect 425610 110898 425846 111134
rect 456330 111218 456566 111454
rect 456330 110898 456566 111134
rect 487050 111218 487286 111454
rect 487050 110898 487286 111134
rect 517770 111218 518006 111454
rect 517770 110898 518006 111134
rect 548490 111218 548726 111454
rect 548490 110898 548726 111134
rect 24146 97538 24382 97774
rect 24466 97538 24702 97774
rect 24146 97218 24382 97454
rect 24466 97218 24702 97454
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 41610 78938 41846 79174
rect 41610 78618 41846 78854
rect 72330 78938 72566 79174
rect 72330 78618 72566 78854
rect 103050 78938 103286 79174
rect 103050 78618 103286 78854
rect 133770 78938 134006 79174
rect 133770 78618 134006 78854
rect 164490 78938 164726 79174
rect 164490 78618 164726 78854
rect 195210 78938 195446 79174
rect 195210 78618 195446 78854
rect 225930 78938 226166 79174
rect 225930 78618 226166 78854
rect 256650 78938 256886 79174
rect 256650 78618 256886 78854
rect 287370 78938 287606 79174
rect 287370 78618 287606 78854
rect 318090 78938 318326 79174
rect 318090 78618 318326 78854
rect 348810 78938 349046 79174
rect 348810 78618 349046 78854
rect 379530 78938 379766 79174
rect 379530 78618 379766 78854
rect 410250 78938 410486 79174
rect 410250 78618 410486 78854
rect 440970 78938 441206 79174
rect 440970 78618 441206 78854
rect 471690 78938 471926 79174
rect 471690 78618 471926 78854
rect 502410 78938 502646 79174
rect 502410 78618 502646 78854
rect 533130 78938 533366 79174
rect 533130 78618 533366 78854
rect 26250 75218 26486 75454
rect 26250 74898 26486 75134
rect 56970 75218 57206 75454
rect 56970 74898 57206 75134
rect 87690 75218 87926 75454
rect 87690 74898 87926 75134
rect 118410 75218 118646 75454
rect 118410 74898 118646 75134
rect 149130 75218 149366 75454
rect 149130 74898 149366 75134
rect 179850 75218 180086 75454
rect 179850 74898 180086 75134
rect 210570 75218 210806 75454
rect 210570 74898 210806 75134
rect 241290 75218 241526 75454
rect 241290 74898 241526 75134
rect 272010 75218 272246 75454
rect 272010 74898 272246 75134
rect 302730 75218 302966 75454
rect 302730 74898 302966 75134
rect 333450 75218 333686 75454
rect 333450 74898 333686 75134
rect 364170 75218 364406 75454
rect 364170 74898 364406 75134
rect 394890 75218 395126 75454
rect 394890 74898 395126 75134
rect 425610 75218 425846 75454
rect 425610 74898 425846 75134
rect 456330 75218 456566 75454
rect 456330 74898 456566 75134
rect 487050 75218 487286 75454
rect 487050 74898 487286 75134
rect 517770 75218 518006 75454
rect 517770 74898 518006 75134
rect 548490 75218 548726 75454
rect 548490 74898 548726 75134
rect 24146 61538 24382 61774
rect 24466 61538 24702 61774
rect 24146 61218 24382 61454
rect 24466 61218 24702 61454
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 41610 42938 41846 43174
rect 41610 42618 41846 42854
rect 72330 42938 72566 43174
rect 72330 42618 72566 42854
rect 103050 42938 103286 43174
rect 103050 42618 103286 42854
rect 133770 42938 134006 43174
rect 133770 42618 134006 42854
rect 164490 42938 164726 43174
rect 164490 42618 164726 42854
rect 195210 42938 195446 43174
rect 195210 42618 195446 42854
rect 225930 42938 226166 43174
rect 225930 42618 226166 42854
rect 256650 42938 256886 43174
rect 256650 42618 256886 42854
rect 287370 42938 287606 43174
rect 287370 42618 287606 42854
rect 318090 42938 318326 43174
rect 318090 42618 318326 42854
rect 348810 42938 349046 43174
rect 348810 42618 349046 42854
rect 379530 42938 379766 43174
rect 379530 42618 379766 42854
rect 410250 42938 410486 43174
rect 410250 42618 410486 42854
rect 440970 42938 441206 43174
rect 440970 42618 441206 42854
rect 471690 42938 471926 43174
rect 471690 42618 471926 42854
rect 502410 42938 502646 43174
rect 502410 42618 502646 42854
rect 533130 42938 533366 43174
rect 533130 42618 533366 42854
rect 26250 39218 26486 39454
rect 26250 38898 26486 39134
rect 56970 39218 57206 39454
rect 56970 38898 57206 39134
rect 87690 39218 87926 39454
rect 87690 38898 87926 39134
rect 118410 39218 118646 39454
rect 118410 38898 118646 39134
rect 149130 39218 149366 39454
rect 149130 38898 149366 39134
rect 179850 39218 180086 39454
rect 179850 38898 180086 39134
rect 210570 39218 210806 39454
rect 210570 38898 210806 39134
rect 241290 39218 241526 39454
rect 241290 38898 241526 39134
rect 272010 39218 272246 39454
rect 272010 38898 272246 39134
rect 302730 39218 302966 39454
rect 302730 38898 302966 39134
rect 333450 39218 333686 39454
rect 333450 38898 333686 39134
rect 364170 39218 364406 39454
rect 364170 38898 364406 39134
rect 394890 39218 395126 39454
rect 394890 38898 395126 39134
rect 425610 39218 425846 39454
rect 425610 38898 425846 39134
rect 456330 39218 456566 39454
rect 456330 38898 456566 39134
rect 487050 39218 487286 39454
rect 487050 38898 487286 39134
rect 517770 39218 518006 39454
rect 517770 38898 518006 39134
rect 548490 39218 548726 39454
rect 548490 38898 548726 39134
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 21649 56662 21885
rect 56746 21649 56982 21885
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 21649 164662 21885
rect 164746 21649 164982 21885
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41610 655174
rect 41846 654938 72330 655174
rect 72566 654938 103050 655174
rect 103286 654938 133770 655174
rect 134006 654938 164490 655174
rect 164726 654938 195210 655174
rect 195446 654938 225930 655174
rect 226166 654938 256650 655174
rect 256886 654938 287370 655174
rect 287606 654938 318090 655174
rect 318326 654938 348810 655174
rect 349046 654938 379530 655174
rect 379766 654938 410250 655174
rect 410486 654938 440970 655174
rect 441206 654938 471690 655174
rect 471926 654938 502410 655174
rect 502646 654938 533130 655174
rect 533366 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41610 654854
rect 41846 654618 72330 654854
rect 72566 654618 103050 654854
rect 103286 654618 133770 654854
rect 134006 654618 164490 654854
rect 164726 654618 195210 654854
rect 195446 654618 225930 654854
rect 226166 654618 256650 654854
rect 256886 654618 287370 654854
rect 287606 654618 318090 654854
rect 318326 654618 348810 654854
rect 349046 654618 379530 654854
rect 379766 654618 410250 654854
rect 410486 654618 440970 654854
rect 441206 654618 471690 654854
rect 471926 654618 502410 654854
rect 502646 654618 533130 654854
rect 533366 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 26250 651454
rect 26486 651218 56970 651454
rect 57206 651218 87690 651454
rect 87926 651218 118410 651454
rect 118646 651218 149130 651454
rect 149366 651218 179850 651454
rect 180086 651218 210570 651454
rect 210806 651218 241290 651454
rect 241526 651218 272010 651454
rect 272246 651218 302730 651454
rect 302966 651218 333450 651454
rect 333686 651218 364170 651454
rect 364406 651218 394890 651454
rect 395126 651218 425610 651454
rect 425846 651218 456330 651454
rect 456566 651218 487050 651454
rect 487286 651218 517770 651454
rect 518006 651218 548490 651454
rect 548726 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 26250 651134
rect 26486 650898 56970 651134
rect 57206 650898 87690 651134
rect 87926 650898 118410 651134
rect 118646 650898 149130 651134
rect 149366 650898 179850 651134
rect 180086 650898 210570 651134
rect 210806 650898 241290 651134
rect 241526 650898 272010 651134
rect 272246 650898 302730 651134
rect 302966 650898 333450 651134
rect 333686 650898 364170 651134
rect 364406 650898 394890 651134
rect 395126 650898 425610 651134
rect 425846 650898 456330 651134
rect 456566 650898 487050 651134
rect 487286 650898 517770 651134
rect 518006 650898 548490 651134
rect 548726 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41610 619174
rect 41846 618938 72330 619174
rect 72566 618938 103050 619174
rect 103286 618938 133770 619174
rect 134006 618938 164490 619174
rect 164726 618938 195210 619174
rect 195446 618938 225930 619174
rect 226166 618938 256650 619174
rect 256886 618938 287370 619174
rect 287606 618938 318090 619174
rect 318326 618938 348810 619174
rect 349046 618938 379530 619174
rect 379766 618938 410250 619174
rect 410486 618938 440970 619174
rect 441206 618938 471690 619174
rect 471926 618938 502410 619174
rect 502646 618938 533130 619174
rect 533366 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41610 618854
rect 41846 618618 72330 618854
rect 72566 618618 103050 618854
rect 103286 618618 133770 618854
rect 134006 618618 164490 618854
rect 164726 618618 195210 618854
rect 195446 618618 225930 618854
rect 226166 618618 256650 618854
rect 256886 618618 287370 618854
rect 287606 618618 318090 618854
rect 318326 618618 348810 618854
rect 349046 618618 379530 618854
rect 379766 618618 410250 618854
rect 410486 618618 440970 618854
rect 441206 618618 471690 618854
rect 471926 618618 502410 618854
rect 502646 618618 533130 618854
rect 533366 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 26250 615454
rect 26486 615218 56970 615454
rect 57206 615218 87690 615454
rect 87926 615218 118410 615454
rect 118646 615218 149130 615454
rect 149366 615218 179850 615454
rect 180086 615218 210570 615454
rect 210806 615218 241290 615454
rect 241526 615218 272010 615454
rect 272246 615218 302730 615454
rect 302966 615218 333450 615454
rect 333686 615218 364170 615454
rect 364406 615218 394890 615454
rect 395126 615218 425610 615454
rect 425846 615218 456330 615454
rect 456566 615218 487050 615454
rect 487286 615218 517770 615454
rect 518006 615218 548490 615454
rect 548726 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 26250 615134
rect 26486 614898 56970 615134
rect 57206 614898 87690 615134
rect 87926 614898 118410 615134
rect 118646 614898 149130 615134
rect 149366 614898 179850 615134
rect 180086 614898 210570 615134
rect 210806 614898 241290 615134
rect 241526 614898 272010 615134
rect 272246 614898 302730 615134
rect 302966 614898 333450 615134
rect 333686 614898 364170 615134
rect 364406 614898 394890 615134
rect 395126 614898 425610 615134
rect 425846 614898 456330 615134
rect 456566 614898 487050 615134
rect 487286 614898 517770 615134
rect 518006 614898 548490 615134
rect 548726 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41610 583174
rect 41846 582938 72330 583174
rect 72566 582938 103050 583174
rect 103286 582938 133770 583174
rect 134006 582938 164490 583174
rect 164726 582938 195210 583174
rect 195446 582938 225930 583174
rect 226166 582938 256650 583174
rect 256886 582938 287370 583174
rect 287606 582938 318090 583174
rect 318326 582938 348810 583174
rect 349046 582938 379530 583174
rect 379766 582938 410250 583174
rect 410486 582938 440970 583174
rect 441206 582938 471690 583174
rect 471926 582938 502410 583174
rect 502646 582938 533130 583174
rect 533366 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41610 582854
rect 41846 582618 72330 582854
rect 72566 582618 103050 582854
rect 103286 582618 133770 582854
rect 134006 582618 164490 582854
rect 164726 582618 195210 582854
rect 195446 582618 225930 582854
rect 226166 582618 256650 582854
rect 256886 582618 287370 582854
rect 287606 582618 318090 582854
rect 318326 582618 348810 582854
rect 349046 582618 379530 582854
rect 379766 582618 410250 582854
rect 410486 582618 440970 582854
rect 441206 582618 471690 582854
rect 471926 582618 502410 582854
rect 502646 582618 533130 582854
rect 533366 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 26250 579454
rect 26486 579218 56970 579454
rect 57206 579218 87690 579454
rect 87926 579218 118410 579454
rect 118646 579218 149130 579454
rect 149366 579218 179850 579454
rect 180086 579218 210570 579454
rect 210806 579218 241290 579454
rect 241526 579218 272010 579454
rect 272246 579218 302730 579454
rect 302966 579218 333450 579454
rect 333686 579218 364170 579454
rect 364406 579218 394890 579454
rect 395126 579218 425610 579454
rect 425846 579218 456330 579454
rect 456566 579218 487050 579454
rect 487286 579218 517770 579454
rect 518006 579218 548490 579454
rect 548726 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 26250 579134
rect 26486 578898 56970 579134
rect 57206 578898 87690 579134
rect 87926 578898 118410 579134
rect 118646 578898 149130 579134
rect 149366 578898 179850 579134
rect 180086 578898 210570 579134
rect 210806 578898 241290 579134
rect 241526 578898 272010 579134
rect 272246 578898 302730 579134
rect 302966 578898 333450 579134
rect 333686 578898 364170 579134
rect 364406 578898 394890 579134
rect 395126 578898 425610 579134
rect 425846 578898 456330 579134
rect 456566 578898 487050 579134
rect 487286 578898 517770 579134
rect 518006 578898 548490 579134
rect 548726 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41610 547174
rect 41846 546938 72330 547174
rect 72566 546938 103050 547174
rect 103286 546938 133770 547174
rect 134006 546938 164490 547174
rect 164726 546938 195210 547174
rect 195446 546938 225930 547174
rect 226166 546938 256650 547174
rect 256886 546938 287370 547174
rect 287606 546938 318090 547174
rect 318326 546938 348810 547174
rect 349046 546938 379530 547174
rect 379766 546938 410250 547174
rect 410486 546938 440970 547174
rect 441206 546938 471690 547174
rect 471926 546938 502410 547174
rect 502646 546938 533130 547174
rect 533366 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41610 546854
rect 41846 546618 72330 546854
rect 72566 546618 103050 546854
rect 103286 546618 133770 546854
rect 134006 546618 164490 546854
rect 164726 546618 195210 546854
rect 195446 546618 225930 546854
rect 226166 546618 256650 546854
rect 256886 546618 287370 546854
rect 287606 546618 318090 546854
rect 318326 546618 348810 546854
rect 349046 546618 379530 546854
rect 379766 546618 410250 546854
rect 410486 546618 440970 546854
rect 441206 546618 471690 546854
rect 471926 546618 502410 546854
rect 502646 546618 533130 546854
rect 533366 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 26250 543454
rect 26486 543218 56970 543454
rect 57206 543218 87690 543454
rect 87926 543218 118410 543454
rect 118646 543218 149130 543454
rect 149366 543218 179850 543454
rect 180086 543218 210570 543454
rect 210806 543218 241290 543454
rect 241526 543218 272010 543454
rect 272246 543218 302730 543454
rect 302966 543218 333450 543454
rect 333686 543218 364170 543454
rect 364406 543218 394890 543454
rect 395126 543218 425610 543454
rect 425846 543218 456330 543454
rect 456566 543218 487050 543454
rect 487286 543218 517770 543454
rect 518006 543218 548490 543454
rect 548726 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 26250 543134
rect 26486 542898 56970 543134
rect 57206 542898 87690 543134
rect 87926 542898 118410 543134
rect 118646 542898 149130 543134
rect 149366 542898 179850 543134
rect 180086 542898 210570 543134
rect 210806 542898 241290 543134
rect 241526 542898 272010 543134
rect 272246 542898 302730 543134
rect 302966 542898 333450 543134
rect 333686 542898 364170 543134
rect 364406 542898 394890 543134
rect 395126 542898 425610 543134
rect 425846 542898 456330 543134
rect 456566 542898 487050 543134
rect 487286 542898 517770 543134
rect 518006 542898 548490 543134
rect 548726 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41610 511174
rect 41846 510938 72330 511174
rect 72566 510938 103050 511174
rect 103286 510938 133770 511174
rect 134006 510938 164490 511174
rect 164726 510938 195210 511174
rect 195446 510938 225930 511174
rect 226166 510938 256650 511174
rect 256886 510938 287370 511174
rect 287606 510938 318090 511174
rect 318326 510938 348810 511174
rect 349046 510938 379530 511174
rect 379766 510938 410250 511174
rect 410486 510938 440970 511174
rect 441206 510938 471690 511174
rect 471926 510938 502410 511174
rect 502646 510938 533130 511174
rect 533366 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41610 510854
rect 41846 510618 72330 510854
rect 72566 510618 103050 510854
rect 103286 510618 133770 510854
rect 134006 510618 164490 510854
rect 164726 510618 195210 510854
rect 195446 510618 225930 510854
rect 226166 510618 256650 510854
rect 256886 510618 287370 510854
rect 287606 510618 318090 510854
rect 318326 510618 348810 510854
rect 349046 510618 379530 510854
rect 379766 510618 410250 510854
rect 410486 510618 440970 510854
rect 441206 510618 471690 510854
rect 471926 510618 502410 510854
rect 502646 510618 533130 510854
rect 533366 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 26250 507454
rect 26486 507218 56970 507454
rect 57206 507218 87690 507454
rect 87926 507218 118410 507454
rect 118646 507218 149130 507454
rect 149366 507218 179850 507454
rect 180086 507218 210570 507454
rect 210806 507218 241290 507454
rect 241526 507218 272010 507454
rect 272246 507218 302730 507454
rect 302966 507218 333450 507454
rect 333686 507218 364170 507454
rect 364406 507218 394890 507454
rect 395126 507218 425610 507454
rect 425846 507218 456330 507454
rect 456566 507218 487050 507454
rect 487286 507218 517770 507454
rect 518006 507218 548490 507454
rect 548726 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 26250 507134
rect 26486 506898 56970 507134
rect 57206 506898 87690 507134
rect 87926 506898 118410 507134
rect 118646 506898 149130 507134
rect 149366 506898 179850 507134
rect 180086 506898 210570 507134
rect 210806 506898 241290 507134
rect 241526 506898 272010 507134
rect 272246 506898 302730 507134
rect 302966 506898 333450 507134
rect 333686 506898 364170 507134
rect 364406 506898 394890 507134
rect 395126 506898 425610 507134
rect 425846 506898 456330 507134
rect 456566 506898 487050 507134
rect 487286 506898 517770 507134
rect 518006 506898 548490 507134
rect 548726 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41610 475174
rect 41846 474938 72330 475174
rect 72566 474938 103050 475174
rect 103286 474938 133770 475174
rect 134006 474938 164490 475174
rect 164726 474938 195210 475174
rect 195446 474938 225930 475174
rect 226166 474938 256650 475174
rect 256886 474938 287370 475174
rect 287606 474938 318090 475174
rect 318326 474938 348810 475174
rect 349046 474938 379530 475174
rect 379766 474938 410250 475174
rect 410486 474938 440970 475174
rect 441206 474938 471690 475174
rect 471926 474938 502410 475174
rect 502646 474938 533130 475174
rect 533366 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41610 474854
rect 41846 474618 72330 474854
rect 72566 474618 103050 474854
rect 103286 474618 133770 474854
rect 134006 474618 164490 474854
rect 164726 474618 195210 474854
rect 195446 474618 225930 474854
rect 226166 474618 256650 474854
rect 256886 474618 287370 474854
rect 287606 474618 318090 474854
rect 318326 474618 348810 474854
rect 349046 474618 379530 474854
rect 379766 474618 410250 474854
rect 410486 474618 440970 474854
rect 441206 474618 471690 474854
rect 471926 474618 502410 474854
rect 502646 474618 533130 474854
rect 533366 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 26250 471454
rect 26486 471218 56970 471454
rect 57206 471218 87690 471454
rect 87926 471218 118410 471454
rect 118646 471218 149130 471454
rect 149366 471218 179850 471454
rect 180086 471218 210570 471454
rect 210806 471218 241290 471454
rect 241526 471218 272010 471454
rect 272246 471218 302730 471454
rect 302966 471218 333450 471454
rect 333686 471218 364170 471454
rect 364406 471218 394890 471454
rect 395126 471218 425610 471454
rect 425846 471218 456330 471454
rect 456566 471218 487050 471454
rect 487286 471218 517770 471454
rect 518006 471218 548490 471454
rect 548726 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 26250 471134
rect 26486 470898 56970 471134
rect 57206 470898 87690 471134
rect 87926 470898 118410 471134
rect 118646 470898 149130 471134
rect 149366 470898 179850 471134
rect 180086 470898 210570 471134
rect 210806 470898 241290 471134
rect 241526 470898 272010 471134
rect 272246 470898 302730 471134
rect 302966 470898 333450 471134
rect 333686 470898 364170 471134
rect 364406 470898 394890 471134
rect 395126 470898 425610 471134
rect 425846 470898 456330 471134
rect 456566 470898 487050 471134
rect 487286 470898 517770 471134
rect 518006 470898 548490 471134
rect 548726 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41610 439174
rect 41846 438938 72330 439174
rect 72566 438938 103050 439174
rect 103286 438938 133770 439174
rect 134006 438938 164490 439174
rect 164726 438938 195210 439174
rect 195446 438938 225930 439174
rect 226166 438938 256650 439174
rect 256886 438938 287370 439174
rect 287606 438938 318090 439174
rect 318326 438938 348810 439174
rect 349046 438938 379530 439174
rect 379766 438938 410250 439174
rect 410486 438938 440970 439174
rect 441206 438938 471690 439174
rect 471926 438938 502410 439174
rect 502646 438938 533130 439174
rect 533366 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41610 438854
rect 41846 438618 72330 438854
rect 72566 438618 103050 438854
rect 103286 438618 133770 438854
rect 134006 438618 164490 438854
rect 164726 438618 195210 438854
rect 195446 438618 225930 438854
rect 226166 438618 256650 438854
rect 256886 438618 287370 438854
rect 287606 438618 318090 438854
rect 318326 438618 348810 438854
rect 349046 438618 379530 438854
rect 379766 438618 410250 438854
rect 410486 438618 440970 438854
rect 441206 438618 471690 438854
rect 471926 438618 502410 438854
rect 502646 438618 533130 438854
rect 533366 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 26250 435454
rect 26486 435218 56970 435454
rect 57206 435218 87690 435454
rect 87926 435218 118410 435454
rect 118646 435218 149130 435454
rect 149366 435218 179850 435454
rect 180086 435218 210570 435454
rect 210806 435218 241290 435454
rect 241526 435218 272010 435454
rect 272246 435218 302730 435454
rect 302966 435218 333450 435454
rect 333686 435218 364170 435454
rect 364406 435218 394890 435454
rect 395126 435218 425610 435454
rect 425846 435218 456330 435454
rect 456566 435218 487050 435454
rect 487286 435218 517770 435454
rect 518006 435218 548490 435454
rect 548726 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 26250 435134
rect 26486 434898 56970 435134
rect 57206 434898 87690 435134
rect 87926 434898 118410 435134
rect 118646 434898 149130 435134
rect 149366 434898 179850 435134
rect 180086 434898 210570 435134
rect 210806 434898 241290 435134
rect 241526 434898 272010 435134
rect 272246 434898 302730 435134
rect 302966 434898 333450 435134
rect 333686 434898 364170 435134
rect 364406 434898 394890 435134
rect 395126 434898 425610 435134
rect 425846 434898 456330 435134
rect 456566 434898 487050 435134
rect 487286 434898 517770 435134
rect 518006 434898 548490 435134
rect 548726 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41610 403174
rect 41846 402938 72330 403174
rect 72566 402938 103050 403174
rect 103286 402938 133770 403174
rect 134006 402938 164490 403174
rect 164726 402938 195210 403174
rect 195446 402938 225930 403174
rect 226166 402938 256650 403174
rect 256886 402938 287370 403174
rect 287606 402938 318090 403174
rect 318326 402938 348810 403174
rect 349046 402938 379530 403174
rect 379766 402938 410250 403174
rect 410486 402938 440970 403174
rect 441206 402938 471690 403174
rect 471926 402938 502410 403174
rect 502646 402938 533130 403174
rect 533366 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41610 402854
rect 41846 402618 72330 402854
rect 72566 402618 103050 402854
rect 103286 402618 133770 402854
rect 134006 402618 164490 402854
rect 164726 402618 195210 402854
rect 195446 402618 225930 402854
rect 226166 402618 256650 402854
rect 256886 402618 287370 402854
rect 287606 402618 318090 402854
rect 318326 402618 348810 402854
rect 349046 402618 379530 402854
rect 379766 402618 410250 402854
rect 410486 402618 440970 402854
rect 441206 402618 471690 402854
rect 471926 402618 502410 402854
rect 502646 402618 533130 402854
rect 533366 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 26250 399454
rect 26486 399218 56970 399454
rect 57206 399218 87690 399454
rect 87926 399218 118410 399454
rect 118646 399218 149130 399454
rect 149366 399218 179850 399454
rect 180086 399218 210570 399454
rect 210806 399218 241290 399454
rect 241526 399218 272010 399454
rect 272246 399218 302730 399454
rect 302966 399218 333450 399454
rect 333686 399218 364170 399454
rect 364406 399218 394890 399454
rect 395126 399218 425610 399454
rect 425846 399218 456330 399454
rect 456566 399218 487050 399454
rect 487286 399218 517770 399454
rect 518006 399218 548490 399454
rect 548726 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 26250 399134
rect 26486 398898 56970 399134
rect 57206 398898 87690 399134
rect 87926 398898 118410 399134
rect 118646 398898 149130 399134
rect 149366 398898 179850 399134
rect 180086 398898 210570 399134
rect 210806 398898 241290 399134
rect 241526 398898 272010 399134
rect 272246 398898 302730 399134
rect 302966 398898 333450 399134
rect 333686 398898 364170 399134
rect 364406 398898 394890 399134
rect 395126 398898 425610 399134
rect 425846 398898 456330 399134
rect 456566 398898 487050 399134
rect 487286 398898 517770 399134
rect 518006 398898 548490 399134
rect 548726 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41610 367174
rect 41846 366938 72330 367174
rect 72566 366938 103050 367174
rect 103286 366938 133770 367174
rect 134006 366938 164490 367174
rect 164726 366938 195210 367174
rect 195446 366938 225930 367174
rect 226166 366938 256650 367174
rect 256886 366938 287370 367174
rect 287606 366938 318090 367174
rect 318326 366938 348810 367174
rect 349046 366938 379530 367174
rect 379766 366938 410250 367174
rect 410486 366938 440970 367174
rect 441206 366938 471690 367174
rect 471926 366938 502410 367174
rect 502646 366938 533130 367174
rect 533366 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41610 366854
rect 41846 366618 72330 366854
rect 72566 366618 103050 366854
rect 103286 366618 133770 366854
rect 134006 366618 164490 366854
rect 164726 366618 195210 366854
rect 195446 366618 225930 366854
rect 226166 366618 256650 366854
rect 256886 366618 287370 366854
rect 287606 366618 318090 366854
rect 318326 366618 348810 366854
rect 349046 366618 379530 366854
rect 379766 366618 410250 366854
rect 410486 366618 440970 366854
rect 441206 366618 471690 366854
rect 471926 366618 502410 366854
rect 502646 366618 533130 366854
rect 533366 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 26250 363454
rect 26486 363218 56970 363454
rect 57206 363218 87690 363454
rect 87926 363218 118410 363454
rect 118646 363218 149130 363454
rect 149366 363218 179850 363454
rect 180086 363218 210570 363454
rect 210806 363218 241290 363454
rect 241526 363218 272010 363454
rect 272246 363218 302730 363454
rect 302966 363218 333450 363454
rect 333686 363218 364170 363454
rect 364406 363218 394890 363454
rect 395126 363218 425610 363454
rect 425846 363218 456330 363454
rect 456566 363218 487050 363454
rect 487286 363218 517770 363454
rect 518006 363218 548490 363454
rect 548726 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 26250 363134
rect 26486 362898 56970 363134
rect 57206 362898 87690 363134
rect 87926 362898 118410 363134
rect 118646 362898 149130 363134
rect 149366 362898 179850 363134
rect 180086 362898 210570 363134
rect 210806 362898 241290 363134
rect 241526 362898 272010 363134
rect 272246 362898 302730 363134
rect 302966 362898 333450 363134
rect 333686 362898 364170 363134
rect 364406 362898 394890 363134
rect 395126 362898 425610 363134
rect 425846 362898 456330 363134
rect 456566 362898 487050 363134
rect 487286 362898 517770 363134
rect 518006 362898 548490 363134
rect 548726 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41610 331174
rect 41846 330938 72330 331174
rect 72566 330938 103050 331174
rect 103286 330938 133770 331174
rect 134006 330938 164490 331174
rect 164726 330938 195210 331174
rect 195446 330938 225930 331174
rect 226166 330938 256650 331174
rect 256886 330938 287370 331174
rect 287606 330938 318090 331174
rect 318326 330938 348810 331174
rect 349046 330938 379530 331174
rect 379766 330938 410250 331174
rect 410486 330938 440970 331174
rect 441206 330938 471690 331174
rect 471926 330938 502410 331174
rect 502646 330938 533130 331174
rect 533366 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41610 330854
rect 41846 330618 72330 330854
rect 72566 330618 103050 330854
rect 103286 330618 133770 330854
rect 134006 330618 164490 330854
rect 164726 330618 195210 330854
rect 195446 330618 225930 330854
rect 226166 330618 256650 330854
rect 256886 330618 287370 330854
rect 287606 330618 318090 330854
rect 318326 330618 348810 330854
rect 349046 330618 379530 330854
rect 379766 330618 410250 330854
rect 410486 330618 440970 330854
rect 441206 330618 471690 330854
rect 471926 330618 502410 330854
rect 502646 330618 533130 330854
rect 533366 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 26250 327454
rect 26486 327218 56970 327454
rect 57206 327218 87690 327454
rect 87926 327218 118410 327454
rect 118646 327218 149130 327454
rect 149366 327218 179850 327454
rect 180086 327218 210570 327454
rect 210806 327218 241290 327454
rect 241526 327218 272010 327454
rect 272246 327218 302730 327454
rect 302966 327218 333450 327454
rect 333686 327218 364170 327454
rect 364406 327218 394890 327454
rect 395126 327218 425610 327454
rect 425846 327218 456330 327454
rect 456566 327218 487050 327454
rect 487286 327218 517770 327454
rect 518006 327218 548490 327454
rect 548726 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 26250 327134
rect 26486 326898 56970 327134
rect 57206 326898 87690 327134
rect 87926 326898 118410 327134
rect 118646 326898 149130 327134
rect 149366 326898 179850 327134
rect 180086 326898 210570 327134
rect 210806 326898 241290 327134
rect 241526 326898 272010 327134
rect 272246 326898 302730 327134
rect 302966 326898 333450 327134
rect 333686 326898 364170 327134
rect 364406 326898 394890 327134
rect 395126 326898 425610 327134
rect 425846 326898 456330 327134
rect 456566 326898 487050 327134
rect 487286 326898 517770 327134
rect 518006 326898 548490 327134
rect 548726 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41610 295174
rect 41846 294938 72330 295174
rect 72566 294938 103050 295174
rect 103286 294938 133770 295174
rect 134006 294938 164490 295174
rect 164726 294938 195210 295174
rect 195446 294938 225930 295174
rect 226166 294938 256650 295174
rect 256886 294938 287370 295174
rect 287606 294938 318090 295174
rect 318326 294938 348810 295174
rect 349046 294938 379530 295174
rect 379766 294938 410250 295174
rect 410486 294938 440970 295174
rect 441206 294938 471690 295174
rect 471926 294938 502410 295174
rect 502646 294938 533130 295174
rect 533366 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41610 294854
rect 41846 294618 72330 294854
rect 72566 294618 103050 294854
rect 103286 294618 133770 294854
rect 134006 294618 164490 294854
rect 164726 294618 195210 294854
rect 195446 294618 225930 294854
rect 226166 294618 256650 294854
rect 256886 294618 287370 294854
rect 287606 294618 318090 294854
rect 318326 294618 348810 294854
rect 349046 294618 379530 294854
rect 379766 294618 410250 294854
rect 410486 294618 440970 294854
rect 441206 294618 471690 294854
rect 471926 294618 502410 294854
rect 502646 294618 533130 294854
rect 533366 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 26250 291454
rect 26486 291218 56970 291454
rect 57206 291218 87690 291454
rect 87926 291218 118410 291454
rect 118646 291218 149130 291454
rect 149366 291218 179850 291454
rect 180086 291218 210570 291454
rect 210806 291218 241290 291454
rect 241526 291218 272010 291454
rect 272246 291218 302730 291454
rect 302966 291218 333450 291454
rect 333686 291218 364170 291454
rect 364406 291218 394890 291454
rect 395126 291218 425610 291454
rect 425846 291218 456330 291454
rect 456566 291218 487050 291454
rect 487286 291218 517770 291454
rect 518006 291218 548490 291454
rect 548726 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 26250 291134
rect 26486 290898 56970 291134
rect 57206 290898 87690 291134
rect 87926 290898 118410 291134
rect 118646 290898 149130 291134
rect 149366 290898 179850 291134
rect 180086 290898 210570 291134
rect 210806 290898 241290 291134
rect 241526 290898 272010 291134
rect 272246 290898 302730 291134
rect 302966 290898 333450 291134
rect 333686 290898 364170 291134
rect 364406 290898 394890 291134
rect 395126 290898 425610 291134
rect 425846 290898 456330 291134
rect 456566 290898 487050 291134
rect 487286 290898 517770 291134
rect 518006 290898 548490 291134
rect 548726 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41610 259174
rect 41846 258938 72330 259174
rect 72566 258938 103050 259174
rect 103286 258938 133770 259174
rect 134006 258938 164490 259174
rect 164726 258938 195210 259174
rect 195446 258938 225930 259174
rect 226166 258938 256650 259174
rect 256886 258938 287370 259174
rect 287606 258938 318090 259174
rect 318326 258938 348810 259174
rect 349046 258938 379530 259174
rect 379766 258938 410250 259174
rect 410486 258938 440970 259174
rect 441206 258938 471690 259174
rect 471926 258938 502410 259174
rect 502646 258938 533130 259174
rect 533366 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41610 258854
rect 41846 258618 72330 258854
rect 72566 258618 103050 258854
rect 103286 258618 133770 258854
rect 134006 258618 164490 258854
rect 164726 258618 195210 258854
rect 195446 258618 225930 258854
rect 226166 258618 256650 258854
rect 256886 258618 287370 258854
rect 287606 258618 318090 258854
rect 318326 258618 348810 258854
rect 349046 258618 379530 258854
rect 379766 258618 410250 258854
rect 410486 258618 440970 258854
rect 441206 258618 471690 258854
rect 471926 258618 502410 258854
rect 502646 258618 533130 258854
rect 533366 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 26250 255454
rect 26486 255218 56970 255454
rect 57206 255218 87690 255454
rect 87926 255218 118410 255454
rect 118646 255218 149130 255454
rect 149366 255218 179850 255454
rect 180086 255218 210570 255454
rect 210806 255218 241290 255454
rect 241526 255218 272010 255454
rect 272246 255218 302730 255454
rect 302966 255218 333450 255454
rect 333686 255218 364170 255454
rect 364406 255218 394890 255454
rect 395126 255218 425610 255454
rect 425846 255218 456330 255454
rect 456566 255218 487050 255454
rect 487286 255218 517770 255454
rect 518006 255218 548490 255454
rect 548726 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 26250 255134
rect 26486 254898 56970 255134
rect 57206 254898 87690 255134
rect 87926 254898 118410 255134
rect 118646 254898 149130 255134
rect 149366 254898 179850 255134
rect 180086 254898 210570 255134
rect 210806 254898 241290 255134
rect 241526 254898 272010 255134
rect 272246 254898 302730 255134
rect 302966 254898 333450 255134
rect 333686 254898 364170 255134
rect 364406 254898 394890 255134
rect 395126 254898 425610 255134
rect 425846 254898 456330 255134
rect 456566 254898 487050 255134
rect 487286 254898 517770 255134
rect 518006 254898 548490 255134
rect 548726 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41610 223174
rect 41846 222938 72330 223174
rect 72566 222938 103050 223174
rect 103286 222938 133770 223174
rect 134006 222938 164490 223174
rect 164726 222938 195210 223174
rect 195446 222938 225930 223174
rect 226166 222938 256650 223174
rect 256886 222938 287370 223174
rect 287606 222938 318090 223174
rect 318326 222938 348810 223174
rect 349046 222938 379530 223174
rect 379766 222938 410250 223174
rect 410486 222938 440970 223174
rect 441206 222938 471690 223174
rect 471926 222938 502410 223174
rect 502646 222938 533130 223174
rect 533366 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41610 222854
rect 41846 222618 72330 222854
rect 72566 222618 103050 222854
rect 103286 222618 133770 222854
rect 134006 222618 164490 222854
rect 164726 222618 195210 222854
rect 195446 222618 225930 222854
rect 226166 222618 256650 222854
rect 256886 222618 287370 222854
rect 287606 222618 318090 222854
rect 318326 222618 348810 222854
rect 349046 222618 379530 222854
rect 379766 222618 410250 222854
rect 410486 222618 440970 222854
rect 441206 222618 471690 222854
rect 471926 222618 502410 222854
rect 502646 222618 533130 222854
rect 533366 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 26250 219454
rect 26486 219218 56970 219454
rect 57206 219218 87690 219454
rect 87926 219218 118410 219454
rect 118646 219218 149130 219454
rect 149366 219218 179850 219454
rect 180086 219218 210570 219454
rect 210806 219218 241290 219454
rect 241526 219218 272010 219454
rect 272246 219218 302730 219454
rect 302966 219218 333450 219454
rect 333686 219218 364170 219454
rect 364406 219218 394890 219454
rect 395126 219218 425610 219454
rect 425846 219218 456330 219454
rect 456566 219218 487050 219454
rect 487286 219218 517770 219454
rect 518006 219218 548490 219454
rect 548726 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 26250 219134
rect 26486 218898 56970 219134
rect 57206 218898 87690 219134
rect 87926 218898 118410 219134
rect 118646 218898 149130 219134
rect 149366 218898 179850 219134
rect 180086 218898 210570 219134
rect 210806 218898 241290 219134
rect 241526 218898 272010 219134
rect 272246 218898 302730 219134
rect 302966 218898 333450 219134
rect 333686 218898 364170 219134
rect 364406 218898 394890 219134
rect 395126 218898 425610 219134
rect 425846 218898 456330 219134
rect 456566 218898 487050 219134
rect 487286 218898 517770 219134
rect 518006 218898 548490 219134
rect 548726 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41610 187174
rect 41846 186938 72330 187174
rect 72566 186938 103050 187174
rect 103286 186938 133770 187174
rect 134006 186938 164490 187174
rect 164726 186938 195210 187174
rect 195446 186938 225930 187174
rect 226166 186938 256650 187174
rect 256886 186938 287370 187174
rect 287606 186938 318090 187174
rect 318326 186938 348810 187174
rect 349046 186938 379530 187174
rect 379766 186938 410250 187174
rect 410486 186938 440970 187174
rect 441206 186938 471690 187174
rect 471926 186938 502410 187174
rect 502646 186938 533130 187174
rect 533366 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41610 186854
rect 41846 186618 72330 186854
rect 72566 186618 103050 186854
rect 103286 186618 133770 186854
rect 134006 186618 164490 186854
rect 164726 186618 195210 186854
rect 195446 186618 225930 186854
rect 226166 186618 256650 186854
rect 256886 186618 287370 186854
rect 287606 186618 318090 186854
rect 318326 186618 348810 186854
rect 349046 186618 379530 186854
rect 379766 186618 410250 186854
rect 410486 186618 440970 186854
rect 441206 186618 471690 186854
rect 471926 186618 502410 186854
rect 502646 186618 533130 186854
rect 533366 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 26250 183454
rect 26486 183218 56970 183454
rect 57206 183218 87690 183454
rect 87926 183218 118410 183454
rect 118646 183218 149130 183454
rect 149366 183218 179850 183454
rect 180086 183218 210570 183454
rect 210806 183218 241290 183454
rect 241526 183218 272010 183454
rect 272246 183218 302730 183454
rect 302966 183218 333450 183454
rect 333686 183218 364170 183454
rect 364406 183218 394890 183454
rect 395126 183218 425610 183454
rect 425846 183218 456330 183454
rect 456566 183218 487050 183454
rect 487286 183218 517770 183454
rect 518006 183218 548490 183454
rect 548726 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 26250 183134
rect 26486 182898 56970 183134
rect 57206 182898 87690 183134
rect 87926 182898 118410 183134
rect 118646 182898 149130 183134
rect 149366 182898 179850 183134
rect 180086 182898 210570 183134
rect 210806 182898 241290 183134
rect 241526 182898 272010 183134
rect 272246 182898 302730 183134
rect 302966 182898 333450 183134
rect 333686 182898 364170 183134
rect 364406 182898 394890 183134
rect 395126 182898 425610 183134
rect 425846 182898 456330 183134
rect 456566 182898 487050 183134
rect 487286 182898 517770 183134
rect 518006 182898 548490 183134
rect 548726 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41610 151174
rect 41846 150938 72330 151174
rect 72566 150938 103050 151174
rect 103286 150938 133770 151174
rect 134006 150938 164490 151174
rect 164726 150938 195210 151174
rect 195446 150938 225930 151174
rect 226166 150938 256650 151174
rect 256886 150938 287370 151174
rect 287606 150938 318090 151174
rect 318326 150938 348810 151174
rect 349046 150938 379530 151174
rect 379766 150938 410250 151174
rect 410486 150938 440970 151174
rect 441206 150938 471690 151174
rect 471926 150938 502410 151174
rect 502646 150938 533130 151174
rect 533366 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41610 150854
rect 41846 150618 72330 150854
rect 72566 150618 103050 150854
rect 103286 150618 133770 150854
rect 134006 150618 164490 150854
rect 164726 150618 195210 150854
rect 195446 150618 225930 150854
rect 226166 150618 256650 150854
rect 256886 150618 287370 150854
rect 287606 150618 318090 150854
rect 318326 150618 348810 150854
rect 349046 150618 379530 150854
rect 379766 150618 410250 150854
rect 410486 150618 440970 150854
rect 441206 150618 471690 150854
rect 471926 150618 502410 150854
rect 502646 150618 533130 150854
rect 533366 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 26250 147454
rect 26486 147218 56970 147454
rect 57206 147218 87690 147454
rect 87926 147218 118410 147454
rect 118646 147218 149130 147454
rect 149366 147218 179850 147454
rect 180086 147218 210570 147454
rect 210806 147218 241290 147454
rect 241526 147218 272010 147454
rect 272246 147218 302730 147454
rect 302966 147218 333450 147454
rect 333686 147218 364170 147454
rect 364406 147218 394890 147454
rect 395126 147218 425610 147454
rect 425846 147218 456330 147454
rect 456566 147218 487050 147454
rect 487286 147218 517770 147454
rect 518006 147218 548490 147454
rect 548726 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 26250 147134
rect 26486 146898 56970 147134
rect 57206 146898 87690 147134
rect 87926 146898 118410 147134
rect 118646 146898 149130 147134
rect 149366 146898 179850 147134
rect 180086 146898 210570 147134
rect 210806 146898 241290 147134
rect 241526 146898 272010 147134
rect 272246 146898 302730 147134
rect 302966 146898 333450 147134
rect 333686 146898 364170 147134
rect 364406 146898 394890 147134
rect 395126 146898 425610 147134
rect 425846 146898 456330 147134
rect 456566 146898 487050 147134
rect 487286 146898 517770 147134
rect 518006 146898 548490 147134
rect 548726 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41610 115174
rect 41846 114938 72330 115174
rect 72566 114938 103050 115174
rect 103286 114938 133770 115174
rect 134006 114938 164490 115174
rect 164726 114938 195210 115174
rect 195446 114938 225930 115174
rect 226166 114938 256650 115174
rect 256886 114938 287370 115174
rect 287606 114938 318090 115174
rect 318326 114938 348810 115174
rect 349046 114938 379530 115174
rect 379766 114938 410250 115174
rect 410486 114938 440970 115174
rect 441206 114938 471690 115174
rect 471926 114938 502410 115174
rect 502646 114938 533130 115174
rect 533366 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41610 114854
rect 41846 114618 72330 114854
rect 72566 114618 103050 114854
rect 103286 114618 133770 114854
rect 134006 114618 164490 114854
rect 164726 114618 195210 114854
rect 195446 114618 225930 114854
rect 226166 114618 256650 114854
rect 256886 114618 287370 114854
rect 287606 114618 318090 114854
rect 318326 114618 348810 114854
rect 349046 114618 379530 114854
rect 379766 114618 410250 114854
rect 410486 114618 440970 114854
rect 441206 114618 471690 114854
rect 471926 114618 502410 114854
rect 502646 114618 533130 114854
rect 533366 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 26250 111454
rect 26486 111218 56970 111454
rect 57206 111218 87690 111454
rect 87926 111218 118410 111454
rect 118646 111218 149130 111454
rect 149366 111218 179850 111454
rect 180086 111218 210570 111454
rect 210806 111218 241290 111454
rect 241526 111218 272010 111454
rect 272246 111218 302730 111454
rect 302966 111218 333450 111454
rect 333686 111218 364170 111454
rect 364406 111218 394890 111454
rect 395126 111218 425610 111454
rect 425846 111218 456330 111454
rect 456566 111218 487050 111454
rect 487286 111218 517770 111454
rect 518006 111218 548490 111454
rect 548726 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 26250 111134
rect 26486 110898 56970 111134
rect 57206 110898 87690 111134
rect 87926 110898 118410 111134
rect 118646 110898 149130 111134
rect 149366 110898 179850 111134
rect 180086 110898 210570 111134
rect 210806 110898 241290 111134
rect 241526 110898 272010 111134
rect 272246 110898 302730 111134
rect 302966 110898 333450 111134
rect 333686 110898 364170 111134
rect 364406 110898 394890 111134
rect 395126 110898 425610 111134
rect 425846 110898 456330 111134
rect 456566 110898 487050 111134
rect 487286 110898 517770 111134
rect 518006 110898 548490 111134
rect 548726 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41610 79174
rect 41846 78938 72330 79174
rect 72566 78938 103050 79174
rect 103286 78938 133770 79174
rect 134006 78938 164490 79174
rect 164726 78938 195210 79174
rect 195446 78938 225930 79174
rect 226166 78938 256650 79174
rect 256886 78938 287370 79174
rect 287606 78938 318090 79174
rect 318326 78938 348810 79174
rect 349046 78938 379530 79174
rect 379766 78938 410250 79174
rect 410486 78938 440970 79174
rect 441206 78938 471690 79174
rect 471926 78938 502410 79174
rect 502646 78938 533130 79174
rect 533366 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41610 78854
rect 41846 78618 72330 78854
rect 72566 78618 103050 78854
rect 103286 78618 133770 78854
rect 134006 78618 164490 78854
rect 164726 78618 195210 78854
rect 195446 78618 225930 78854
rect 226166 78618 256650 78854
rect 256886 78618 287370 78854
rect 287606 78618 318090 78854
rect 318326 78618 348810 78854
rect 349046 78618 379530 78854
rect 379766 78618 410250 78854
rect 410486 78618 440970 78854
rect 441206 78618 471690 78854
rect 471926 78618 502410 78854
rect 502646 78618 533130 78854
rect 533366 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 26250 75454
rect 26486 75218 56970 75454
rect 57206 75218 87690 75454
rect 87926 75218 118410 75454
rect 118646 75218 149130 75454
rect 149366 75218 179850 75454
rect 180086 75218 210570 75454
rect 210806 75218 241290 75454
rect 241526 75218 272010 75454
rect 272246 75218 302730 75454
rect 302966 75218 333450 75454
rect 333686 75218 364170 75454
rect 364406 75218 394890 75454
rect 395126 75218 425610 75454
rect 425846 75218 456330 75454
rect 456566 75218 487050 75454
rect 487286 75218 517770 75454
rect 518006 75218 548490 75454
rect 548726 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 26250 75134
rect 26486 74898 56970 75134
rect 57206 74898 87690 75134
rect 87926 74898 118410 75134
rect 118646 74898 149130 75134
rect 149366 74898 179850 75134
rect 180086 74898 210570 75134
rect 210806 74898 241290 75134
rect 241526 74898 272010 75134
rect 272246 74898 302730 75134
rect 302966 74898 333450 75134
rect 333686 74898 364170 75134
rect 364406 74898 394890 75134
rect 395126 74898 425610 75134
rect 425846 74898 456330 75134
rect 456566 74898 487050 75134
rect 487286 74898 517770 75134
rect 518006 74898 548490 75134
rect 548726 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41610 43174
rect 41846 42938 72330 43174
rect 72566 42938 103050 43174
rect 103286 42938 133770 43174
rect 134006 42938 164490 43174
rect 164726 42938 195210 43174
rect 195446 42938 225930 43174
rect 226166 42938 256650 43174
rect 256886 42938 287370 43174
rect 287606 42938 318090 43174
rect 318326 42938 348810 43174
rect 349046 42938 379530 43174
rect 379766 42938 410250 43174
rect 410486 42938 440970 43174
rect 441206 42938 471690 43174
rect 471926 42938 502410 43174
rect 502646 42938 533130 43174
rect 533366 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41610 42854
rect 41846 42618 72330 42854
rect 72566 42618 103050 42854
rect 103286 42618 133770 42854
rect 134006 42618 164490 42854
rect 164726 42618 195210 42854
rect 195446 42618 225930 42854
rect 226166 42618 256650 42854
rect 256886 42618 287370 42854
rect 287606 42618 318090 42854
rect 318326 42618 348810 42854
rect 349046 42618 379530 42854
rect 379766 42618 410250 42854
rect 410486 42618 440970 42854
rect 441206 42618 471690 42854
rect 471926 42618 502410 42854
rect 502646 42618 533130 42854
rect 533366 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 26250 39454
rect 26486 39218 56970 39454
rect 57206 39218 87690 39454
rect 87926 39218 118410 39454
rect 118646 39218 149130 39454
rect 149366 39218 179850 39454
rect 180086 39218 210570 39454
rect 210806 39218 241290 39454
rect 241526 39218 272010 39454
rect 272246 39218 302730 39454
rect 302966 39218 333450 39454
rect 333686 39218 364170 39454
rect 364406 39218 394890 39454
rect 395126 39218 425610 39454
rect 425846 39218 456330 39454
rect 456566 39218 487050 39454
rect 487286 39218 517770 39454
rect 518006 39218 548490 39454
rect 548726 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 26250 39134
rect 26486 38898 56970 39134
rect 57206 38898 87690 39134
rect 87926 38898 118410 39134
rect 118646 38898 149130 39134
rect 149366 38898 179850 39134
rect 180086 38898 210570 39134
rect 210806 38898 241290 39134
rect 241526 38898 272010 39134
rect 272246 38898 302730 39134
rect 302966 38898 333450 39134
rect 333686 38898 364170 39134
rect 364406 38898 394890 39134
rect 395126 38898 425610 39134
rect 425846 38898 456330 39134
rect 456566 38898 487050 39134
rect 487286 38898 517770 39134
rect 518006 38898 548490 39134
rect 548726 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21885 92426 22054
rect 20982 21818 56426 21885
rect -8726 21734 56426 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21649 56426 21734
rect 56662 21649 56746 21885
rect 56982 21818 92426 21885
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21885 200426 22054
rect 128982 21818 164426 21885
rect 56982 21734 164426 21818
rect 56982 21649 92426 21734
rect 20982 21498 92426 21649
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21649 164426 21734
rect 164662 21649 164746 21885
rect 164982 21818 200426 21885
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect 164982 21734 592650 21818
rect 164982 21649 200426 21734
rect 128982 21498 200426 21649
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use WrapperBlock_noparam  mprj
timestamp 0
transform 1 0 22000 0 1 22000
box 0 0 540000 660000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 681449 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 681449 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 681449 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 681449 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 681449 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 681449 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 681449 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 681449 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 681449 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 681449 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 681449 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 681449 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 681449 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 681449 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 22287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 681449 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 681449 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 681449 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 681449 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 681449 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 681449 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 22068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 681804 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 681449 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 681449 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 22068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 681804 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 681449 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 681449 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 22068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 681804 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 681449 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 681449 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 22287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 681449 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 22287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 22068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 22068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 22287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 22068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 681804 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 681449 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 681449 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 681449 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 681449 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 681449 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 681449 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 681449 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 681449 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 681449 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 681449 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 681449 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 681449 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 681449 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 22287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 681449 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 681449 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 681449 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 681449 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 681449 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 681449 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 681449 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 681449 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 681449 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 681449 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 681449 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 681449 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 681449 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 681449 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 681449 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 22287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 681449 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
