VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO VectorRegFile
  CLASS BLOCK ;
  FOREIGN VectorRegFile ;
  ORIGIN 0.000 0.000 ;
  SIZE 1221.615 BY 929.690 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END clk
  PIN rAddr1_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END rAddr1_1[0]
  PIN rAddr1_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END rAddr1_1[1]
  PIN rAddr1_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 925.690 618.610 929.690 ;
    END
  END rAddr1_1[2]
  PIN rAddr1_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 911.240 1221.615 911.840 ;
    END
  END rAddr1_1[3]
  PIN rAddr1_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END rAddr1_1[4]
  PIN rAddr1_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 925.690 1108.050 929.690 ;
    END
  END rAddr1_2[0]
  PIN rAddr1_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END rAddr1_2[1]
  PIN rAddr1_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 925.690 325.590 929.690 ;
    END
  END rAddr1_2[2]
  PIN rAddr1_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END rAddr1_2[3]
  PIN rAddr1_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 925.690 1043.650 929.690 ;
    END
  END rAddr1_2[4]
  PIN rAddr2_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 258.440 1221.615 259.040 ;
    END
  END rAddr2_1[0]
  PIN rAddr2_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 925.690 1075.850 929.690 ;
    END
  END rAddr2_1[1]
  PIN rAddr2_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END rAddr2_1[2]
  PIN rAddr2_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END rAddr2_1[3]
  PIN rAddr2_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 925.690 586.410 929.690 ;
    END
  END rAddr2_1[4]
  PIN rAddr2_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 224.440 1221.615 225.040 ;
    END
  END rAddr2_2[0]
  PIN rAddr2_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 925.690 650.810 929.690 ;
    END
  END rAddr2_2[1]
  PIN rAddr2_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 635.840 1221.615 636.440 ;
    END
  END rAddr2_2[2]
  PIN rAddr2_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END rAddr2_2[3]
  PIN rAddr2_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 465.840 1221.615 466.440 ;
    END
  END rAddr2_2[4]
  PIN rData1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 428.440 1221.615 429.040 ;
    END
  END rData1[0]
  PIN rData1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 925.690 389.990 929.690 ;
    END
  END rData1[10]
  PIN rData1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END rData1[11]
  PIN rData1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END rData1[12]
  PIN rData1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 499.840 1221.615 500.440 ;
    END
  END rData1[13]
  PIN rData1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END rData1[14]
  PIN rData1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END rData1[15]
  PIN rData1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END rData1[16]
  PIN rData1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 601.840 1221.615 602.440 ;
    END
  END rData1[17]
  PIN rData1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 925.690 815.030 929.690 ;
    END
  END rData1[18]
  PIN rData1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END rData1[19]
  PIN rData1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 925.690 257.970 929.690 ;
    END
  END rData1[1]
  PIN rData1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 153.040 1221.615 153.640 ;
    END
  END rData1[20]
  PIN rData1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 925.690 129.170 929.690 ;
    END
  END rData1[21]
  PIN rData1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END rData1[22]
  PIN rData1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 925.690 1172.450 929.690 ;
    END
  END rData1[23]
  PIN rData1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END rData1[24]
  PIN rData1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END rData1[25]
  PIN rData1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END rData1[26]
  PIN rData1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END rData1[27]
  PIN rData1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END rData1[28]
  PIN rData1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 51.040 1221.615 51.640 ;
    END
  END rData1[29]
  PIN rData1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 925.690 747.410 929.690 ;
    END
  END rData1[2]
  PIN rData1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END rData1[30]
  PIN rData1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 925.690 911.630 929.690 ;
    END
  END rData1[31]
  PIN rData1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END rData1[3]
  PIN rData1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 925.690 1204.650 929.690 ;
    END
  END rData1[4]
  PIN rData1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 925.690 454.390 929.690 ;
    END
  END rData1[5]
  PIN rData1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END rData1[6]
  PIN rData1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 669.840 1221.615 670.440 ;
    END
  END rData1[7]
  PIN rData1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END rData1[8]
  PIN rData1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 925.690 715.210 929.690 ;
    END
  END rData1[9]
  PIN rData2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 925.690 518.790 929.690 ;
    END
  END rData2[0]
  PIN rData2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END rData2[10]
  PIN rData2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 877.240 1221.615 877.840 ;
    END
  END rData2[11]
  PIN rData2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END rData2[12]
  PIN rData2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END rData2[13]
  PIN rData2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 925.690 422.190 929.690 ;
    END
  END rData2[14]
  PIN rData2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END rData2[15]
  PIN rData2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 809.240 1221.615 809.840 ;
    END
  END rData2[16]
  PIN rData2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 925.690 225.770 929.690 ;
    END
  END rData2[17]
  PIN rData2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 741.240 1221.615 741.840 ;
    END
  END rData2[18]
  PIN rData2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 925.690 293.390 929.690 ;
    END
  END rData2[19]
  PIN rData2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 925.690 554.210 929.690 ;
    END
  END rData2[1]
  PIN rData2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 925.690 879.430 929.690 ;
    END
  END rData2[20]
  PIN rData2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END rData2[21]
  PIN rData2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 292.440 1221.615 293.040 ;
    END
  END rData2[22]
  PIN rData2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 119.040 1221.615 119.640 ;
    END
  END rData2[23]
  PIN rData2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END rData2[24]
  PIN rData2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END rData2[25]
  PIN rData2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END rData2[26]
  PIN rData2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 190.440 1221.615 191.040 ;
    END
  END rData2[27]
  PIN rData2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END rData2[28]
  PIN rData2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END rData2[29]
  PIN rData2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END rData2[2]
  PIN rData2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END rData2[30]
  PIN rData2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END rData2[31]
  PIN rData2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 843.240 1221.615 843.840 ;
    END
  END rData2[3]
  PIN rData2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END rData2[4]
  PIN rData2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END rData2[5]
  PIN rData2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END rData2[6]
  PIN rData2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END rData2[7]
  PIN rData2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 925.690 683.010 929.690 ;
    END
  END rData2[8]
  PIN rData2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END rData2[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 916.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 916.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 916.880 ;
    END
  END vssd1
  PIN wAddr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END wAddr1[0]
  PIN wAddr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END wAddr1[1]
  PIN wAddr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 567.840 1221.615 568.440 ;
    END
  END wAddr1[2]
  PIN wAddr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 326.440 1221.615 327.040 ;
    END
  END wAddr1[3]
  PIN wAddr1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END wAddr1[4]
  PIN wAddr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END wAddr2[0]
  PIN wAddr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 85.040 1221.615 85.640 ;
    END
  END wAddr2[1]
  PIN wAddr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END wAddr2[2]
  PIN wAddr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 394.440 1221.615 395.040 ;
    END
  END wAddr2[3]
  PIN wAddr2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 707.240 1221.615 707.840 ;
    END
  END wAddr2[4]
  PIN wData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END wData[0]
  PIN wData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 775.240 1221.615 775.840 ;
    END
  END wData[10]
  PIN wData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 925.690 64.770 929.690 ;
    END
  END wData[11]
  PIN wData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END wData[12]
  PIN wData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END wData[13]
  PIN wData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wData[14]
  PIN wData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END wData[15]
  PIN wData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 925.690 161.370 929.690 ;
    END
  END wData[16]
  PIN wData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 925.690 486.590 929.690 ;
    END
  END wData[17]
  PIN wData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 925.690 847.230 929.690 ;
    END
  END wData[18]
  PIN wData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END wData[19]
  PIN wData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END wData[1]
  PIN wData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wData[20]
  PIN wData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 925.690 1011.450 929.690 ;
    END
  END wData[21]
  PIN wData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 925.690 782.830 929.690 ;
    END
  END wData[22]
  PIN wData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END wData[23]
  PIN wData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 925.690 1140.250 929.690 ;
    END
  END wData[24]
  PIN wData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 17.040 1221.615 17.640 ;
    END
  END wData[25]
  PIN wData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 925.690 96.970 929.690 ;
    END
  END wData[26]
  PIN wData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END wData[27]
  PIN wData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wData[28]
  PIN wData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END wData[29]
  PIN wData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END wData[2]
  PIN wData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 533.840 1221.615 534.440 ;
    END
  END wData[30]
  PIN wData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END wData[31]
  PIN wData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 925.690 976.030 929.690 ;
    END
  END wData[3]
  PIN wData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 925.690 943.830 929.690 ;
    END
  END wData[4]
  PIN wData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 925.690 193.570 929.690 ;
    END
  END wData[5]
  PIN wData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 925.690 357.790 929.690 ;
    END
  END wData[6]
  PIN wData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END wData[7]
  PIN wData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END wData[8]
  PIN wData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 925.690 29.350 929.690 ;
    END
  END wData[9]
  PIN wEnable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1217.615 360.440 1221.615 361.040 ;
    END
  END wEnable
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1215.780 916.725 ;
      LAYER met1 ;
        RECT 0.070 4.460 1217.090 925.440 ;
      LAYER met2 ;
        RECT 0.100 925.410 28.790 928.725 ;
        RECT 29.630 925.410 64.210 928.725 ;
        RECT 65.050 925.410 96.410 928.725 ;
        RECT 97.250 925.410 128.610 928.725 ;
        RECT 129.450 925.410 160.810 928.725 ;
        RECT 161.650 925.410 193.010 928.725 ;
        RECT 193.850 925.410 225.210 928.725 ;
        RECT 226.050 925.410 257.410 928.725 ;
        RECT 258.250 925.410 292.830 928.725 ;
        RECT 293.670 925.410 325.030 928.725 ;
        RECT 325.870 925.410 357.230 928.725 ;
        RECT 358.070 925.410 389.430 928.725 ;
        RECT 390.270 925.410 421.630 928.725 ;
        RECT 422.470 925.410 453.830 928.725 ;
        RECT 454.670 925.410 486.030 928.725 ;
        RECT 486.870 925.410 518.230 928.725 ;
        RECT 519.070 925.410 553.650 928.725 ;
        RECT 554.490 925.410 585.850 928.725 ;
        RECT 586.690 925.410 618.050 928.725 ;
        RECT 618.890 925.410 650.250 928.725 ;
        RECT 651.090 925.410 682.450 928.725 ;
        RECT 683.290 925.410 714.650 928.725 ;
        RECT 715.490 925.410 746.850 928.725 ;
        RECT 747.690 925.410 782.270 928.725 ;
        RECT 783.110 925.410 814.470 928.725 ;
        RECT 815.310 925.410 846.670 928.725 ;
        RECT 847.510 925.410 878.870 928.725 ;
        RECT 879.710 925.410 911.070 928.725 ;
        RECT 911.910 925.410 943.270 928.725 ;
        RECT 944.110 925.410 975.470 928.725 ;
        RECT 976.310 925.410 1010.890 928.725 ;
        RECT 1011.730 925.410 1043.090 928.725 ;
        RECT 1043.930 925.410 1075.290 928.725 ;
        RECT 1076.130 925.410 1107.490 928.725 ;
        RECT 1108.330 925.410 1139.690 928.725 ;
        RECT 1140.530 925.410 1171.890 928.725 ;
        RECT 1172.730 925.410 1204.090 928.725 ;
        RECT 1204.930 925.410 1217.070 928.725 ;
        RECT 0.100 4.280 1217.070 925.410 ;
        RECT 0.650 3.670 32.010 4.280 ;
        RECT 32.850 3.670 64.210 4.280 ;
        RECT 65.050 3.670 96.410 4.280 ;
        RECT 97.250 3.670 128.610 4.280 ;
        RECT 129.450 3.670 160.810 4.280 ;
        RECT 161.650 3.670 193.010 4.280 ;
        RECT 193.850 3.670 225.210 4.280 ;
        RECT 226.050 3.670 260.630 4.280 ;
        RECT 261.470 3.670 292.830 4.280 ;
        RECT 293.670 3.670 325.030 4.280 ;
        RECT 325.870 3.670 357.230 4.280 ;
        RECT 358.070 3.670 389.430 4.280 ;
        RECT 390.270 3.670 421.630 4.280 ;
        RECT 422.470 3.670 453.830 4.280 ;
        RECT 454.670 3.670 489.250 4.280 ;
        RECT 490.090 3.670 521.450 4.280 ;
        RECT 522.290 3.670 553.650 4.280 ;
        RECT 554.490 3.670 585.850 4.280 ;
        RECT 586.690 3.670 618.050 4.280 ;
        RECT 618.890 3.670 650.250 4.280 ;
        RECT 651.090 3.670 682.450 4.280 ;
        RECT 683.290 3.670 717.870 4.280 ;
        RECT 718.710 3.670 750.070 4.280 ;
        RECT 750.910 3.670 782.270 4.280 ;
        RECT 783.110 3.670 814.470 4.280 ;
        RECT 815.310 3.670 846.670 4.280 ;
        RECT 847.510 3.670 878.870 4.280 ;
        RECT 879.710 3.670 911.070 4.280 ;
        RECT 911.910 3.670 946.490 4.280 ;
        RECT 947.330 3.670 978.690 4.280 ;
        RECT 979.530 3.670 1010.890 4.280 ;
        RECT 1011.730 3.670 1043.090 4.280 ;
        RECT 1043.930 3.670 1075.290 4.280 ;
        RECT 1076.130 3.670 1107.490 4.280 ;
        RECT 1108.330 3.670 1139.690 4.280 ;
        RECT 1140.530 3.670 1175.110 4.280 ;
        RECT 1175.950 3.670 1207.310 4.280 ;
        RECT 1208.150 3.670 1217.070 4.280 ;
      LAYER met3 ;
        RECT 4.400 927.840 1217.615 928.705 ;
        RECT 4.000 912.240 1217.615 927.840 ;
        RECT 4.000 910.840 1217.215 912.240 ;
        RECT 4.000 895.240 1217.615 910.840 ;
        RECT 4.400 893.840 1217.615 895.240 ;
        RECT 4.000 878.240 1217.615 893.840 ;
        RECT 4.000 876.840 1217.215 878.240 ;
        RECT 4.000 861.240 1217.615 876.840 ;
        RECT 4.400 859.840 1217.615 861.240 ;
        RECT 4.000 844.240 1217.615 859.840 ;
        RECT 4.000 842.840 1217.215 844.240 ;
        RECT 4.000 827.240 1217.615 842.840 ;
        RECT 4.400 825.840 1217.615 827.240 ;
        RECT 4.000 810.240 1217.615 825.840 ;
        RECT 4.000 808.840 1217.215 810.240 ;
        RECT 4.000 793.240 1217.615 808.840 ;
        RECT 4.400 791.840 1217.615 793.240 ;
        RECT 4.000 776.240 1217.615 791.840 ;
        RECT 4.000 774.840 1217.215 776.240 ;
        RECT 4.000 759.240 1217.615 774.840 ;
        RECT 4.400 757.840 1217.615 759.240 ;
        RECT 4.000 742.240 1217.615 757.840 ;
        RECT 4.000 740.840 1217.215 742.240 ;
        RECT 4.000 721.840 1217.615 740.840 ;
        RECT 4.400 720.440 1217.615 721.840 ;
        RECT 4.000 708.240 1217.615 720.440 ;
        RECT 4.000 706.840 1217.215 708.240 ;
        RECT 4.000 687.840 1217.615 706.840 ;
        RECT 4.400 686.440 1217.615 687.840 ;
        RECT 4.000 670.840 1217.615 686.440 ;
        RECT 4.000 669.440 1217.215 670.840 ;
        RECT 4.000 653.840 1217.615 669.440 ;
        RECT 4.400 652.440 1217.615 653.840 ;
        RECT 4.000 636.840 1217.615 652.440 ;
        RECT 4.000 635.440 1217.215 636.840 ;
        RECT 4.000 619.840 1217.615 635.440 ;
        RECT 4.400 618.440 1217.615 619.840 ;
        RECT 4.000 602.840 1217.615 618.440 ;
        RECT 4.000 601.440 1217.215 602.840 ;
        RECT 4.000 585.840 1217.615 601.440 ;
        RECT 4.400 584.440 1217.615 585.840 ;
        RECT 4.000 568.840 1217.615 584.440 ;
        RECT 4.000 567.440 1217.215 568.840 ;
        RECT 4.000 551.840 1217.615 567.440 ;
        RECT 4.400 550.440 1217.615 551.840 ;
        RECT 4.000 534.840 1217.615 550.440 ;
        RECT 4.000 533.440 1217.215 534.840 ;
        RECT 4.000 517.840 1217.615 533.440 ;
        RECT 4.400 516.440 1217.615 517.840 ;
        RECT 4.000 500.840 1217.615 516.440 ;
        RECT 4.000 499.440 1217.215 500.840 ;
        RECT 4.000 480.440 1217.615 499.440 ;
        RECT 4.400 479.040 1217.615 480.440 ;
        RECT 4.000 466.840 1217.615 479.040 ;
        RECT 4.000 465.440 1217.215 466.840 ;
        RECT 4.000 446.440 1217.615 465.440 ;
        RECT 4.400 445.040 1217.615 446.440 ;
        RECT 4.000 429.440 1217.615 445.040 ;
        RECT 4.000 428.040 1217.215 429.440 ;
        RECT 4.000 412.440 1217.615 428.040 ;
        RECT 4.400 411.040 1217.615 412.440 ;
        RECT 4.000 395.440 1217.615 411.040 ;
        RECT 4.000 394.040 1217.215 395.440 ;
        RECT 4.000 378.440 1217.615 394.040 ;
        RECT 4.400 377.040 1217.615 378.440 ;
        RECT 4.000 361.440 1217.615 377.040 ;
        RECT 4.000 360.040 1217.215 361.440 ;
        RECT 4.000 344.440 1217.615 360.040 ;
        RECT 4.400 343.040 1217.615 344.440 ;
        RECT 4.000 327.440 1217.615 343.040 ;
        RECT 4.000 326.040 1217.215 327.440 ;
        RECT 4.000 310.440 1217.615 326.040 ;
        RECT 4.400 309.040 1217.615 310.440 ;
        RECT 4.000 293.440 1217.615 309.040 ;
        RECT 4.000 292.040 1217.215 293.440 ;
        RECT 4.000 276.440 1217.615 292.040 ;
        RECT 4.400 275.040 1217.615 276.440 ;
        RECT 4.000 259.440 1217.615 275.040 ;
        RECT 4.000 258.040 1217.215 259.440 ;
        RECT 4.000 239.040 1217.615 258.040 ;
        RECT 4.400 237.640 1217.615 239.040 ;
        RECT 4.000 225.440 1217.615 237.640 ;
        RECT 4.000 224.040 1217.215 225.440 ;
        RECT 4.000 205.040 1217.615 224.040 ;
        RECT 4.400 203.640 1217.615 205.040 ;
        RECT 4.000 191.440 1217.615 203.640 ;
        RECT 4.000 190.040 1217.215 191.440 ;
        RECT 4.000 171.040 1217.615 190.040 ;
        RECT 4.400 169.640 1217.615 171.040 ;
        RECT 4.000 154.040 1217.615 169.640 ;
        RECT 4.000 152.640 1217.215 154.040 ;
        RECT 4.000 137.040 1217.615 152.640 ;
        RECT 4.400 135.640 1217.615 137.040 ;
        RECT 4.000 120.040 1217.615 135.640 ;
        RECT 4.000 118.640 1217.215 120.040 ;
        RECT 4.000 103.040 1217.615 118.640 ;
        RECT 4.400 101.640 1217.615 103.040 ;
        RECT 4.000 86.040 1217.615 101.640 ;
        RECT 4.000 84.640 1217.215 86.040 ;
        RECT 4.000 69.040 1217.615 84.640 ;
        RECT 4.400 67.640 1217.615 69.040 ;
        RECT 4.000 52.040 1217.615 67.640 ;
        RECT 4.000 50.640 1217.215 52.040 ;
        RECT 4.000 35.040 1217.615 50.640 ;
        RECT 4.400 33.640 1217.615 35.040 ;
        RECT 4.000 18.040 1217.615 33.640 ;
        RECT 4.000 16.640 1217.215 18.040 ;
        RECT 4.000 7.655 1217.615 16.640 ;
      LAYER met4 ;
        RECT 24.215 10.240 97.440 915.785 ;
        RECT 99.840 10.240 174.240 915.785 ;
        RECT 176.640 10.240 251.040 915.785 ;
        RECT 253.440 10.240 327.840 915.785 ;
        RECT 330.240 10.240 404.640 915.785 ;
        RECT 407.040 10.240 481.440 915.785 ;
        RECT 483.840 10.240 558.240 915.785 ;
        RECT 560.640 10.240 635.040 915.785 ;
        RECT 637.440 10.240 711.840 915.785 ;
        RECT 714.240 10.240 788.640 915.785 ;
        RECT 791.040 10.240 865.440 915.785 ;
        RECT 867.840 10.240 942.240 915.785 ;
        RECT 944.640 10.240 1019.040 915.785 ;
        RECT 1021.440 10.240 1095.840 915.785 ;
        RECT 1098.240 10.240 1172.640 915.785 ;
        RECT 1175.040 10.240 1197.545 915.785 ;
        RECT 24.215 7.655 1197.545 10.240 ;
  END
END VectorRegFile
END LIBRARY

