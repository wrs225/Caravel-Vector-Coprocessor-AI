// This is the unpowered netlist.
module Scalar_Register_File (clk,
    reset,
    write_enable,
    read_address,
    read_data,
    write_address,
    write_data);
 input clk;
 input reset;
 input write_enable;
 input [4:0] read_address;
 output [31:0] read_data;
 input [4:0] write_address;
 input [31:0] write_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \srfp.register_file[0][0] ;
 wire \srfp.register_file[0][10] ;
 wire \srfp.register_file[0][11] ;
 wire \srfp.register_file[0][12] ;
 wire \srfp.register_file[0][13] ;
 wire \srfp.register_file[0][14] ;
 wire \srfp.register_file[0][15] ;
 wire \srfp.register_file[0][16] ;
 wire \srfp.register_file[0][17] ;
 wire \srfp.register_file[0][18] ;
 wire \srfp.register_file[0][19] ;
 wire \srfp.register_file[0][1] ;
 wire \srfp.register_file[0][20] ;
 wire \srfp.register_file[0][21] ;
 wire \srfp.register_file[0][22] ;
 wire \srfp.register_file[0][23] ;
 wire \srfp.register_file[0][24] ;
 wire \srfp.register_file[0][25] ;
 wire \srfp.register_file[0][26] ;
 wire \srfp.register_file[0][27] ;
 wire \srfp.register_file[0][28] ;
 wire \srfp.register_file[0][29] ;
 wire \srfp.register_file[0][2] ;
 wire \srfp.register_file[0][30] ;
 wire \srfp.register_file[0][31] ;
 wire \srfp.register_file[0][3] ;
 wire \srfp.register_file[0][4] ;
 wire \srfp.register_file[0][5] ;
 wire \srfp.register_file[0][6] ;
 wire \srfp.register_file[0][7] ;
 wire \srfp.register_file[0][8] ;
 wire \srfp.register_file[0][9] ;
 wire \srfp.register_file[1][0] ;
 wire \srfp.register_file[1][10] ;
 wire \srfp.register_file[1][11] ;
 wire \srfp.register_file[1][12] ;
 wire \srfp.register_file[1][13] ;
 wire \srfp.register_file[1][14] ;
 wire \srfp.register_file[1][15] ;
 wire \srfp.register_file[1][16] ;
 wire \srfp.register_file[1][17] ;
 wire \srfp.register_file[1][18] ;
 wire \srfp.register_file[1][19] ;
 wire \srfp.register_file[1][1] ;
 wire \srfp.register_file[1][20] ;
 wire \srfp.register_file[1][21] ;
 wire \srfp.register_file[1][22] ;
 wire \srfp.register_file[1][23] ;
 wire \srfp.register_file[1][24] ;
 wire \srfp.register_file[1][25] ;
 wire \srfp.register_file[1][26] ;
 wire \srfp.register_file[1][27] ;
 wire \srfp.register_file[1][28] ;
 wire \srfp.register_file[1][29] ;
 wire \srfp.register_file[1][2] ;
 wire \srfp.register_file[1][30] ;
 wire \srfp.register_file[1][31] ;
 wire \srfp.register_file[1][3] ;
 wire \srfp.register_file[1][4] ;
 wire \srfp.register_file[1][5] ;
 wire \srfp.register_file[1][6] ;
 wire \srfp.register_file[1][7] ;
 wire \srfp.register_file[1][8] ;
 wire \srfp.register_file[1][9] ;
 wire \srfp.register_file[2][0] ;
 wire \srfp.register_file[2][10] ;
 wire \srfp.register_file[2][11] ;
 wire \srfp.register_file[2][12] ;
 wire \srfp.register_file[2][13] ;
 wire \srfp.register_file[2][14] ;
 wire \srfp.register_file[2][15] ;
 wire \srfp.register_file[2][16] ;
 wire \srfp.register_file[2][17] ;
 wire \srfp.register_file[2][18] ;
 wire \srfp.register_file[2][19] ;
 wire \srfp.register_file[2][1] ;
 wire \srfp.register_file[2][20] ;
 wire \srfp.register_file[2][21] ;
 wire \srfp.register_file[2][22] ;
 wire \srfp.register_file[2][23] ;
 wire \srfp.register_file[2][24] ;
 wire \srfp.register_file[2][25] ;
 wire \srfp.register_file[2][26] ;
 wire \srfp.register_file[2][27] ;
 wire \srfp.register_file[2][28] ;
 wire \srfp.register_file[2][29] ;
 wire \srfp.register_file[2][2] ;
 wire \srfp.register_file[2][30] ;
 wire \srfp.register_file[2][31] ;
 wire \srfp.register_file[2][3] ;
 wire \srfp.register_file[2][4] ;
 wire \srfp.register_file[2][5] ;
 wire \srfp.register_file[2][6] ;
 wire \srfp.register_file[2][7] ;
 wire \srfp.register_file[2][8] ;
 wire \srfp.register_file[2][9] ;
 wire \srfp.register_file[3][0] ;
 wire \srfp.register_file[3][10] ;
 wire \srfp.register_file[3][11] ;
 wire \srfp.register_file[3][12] ;
 wire \srfp.register_file[3][13] ;
 wire \srfp.register_file[3][14] ;
 wire \srfp.register_file[3][15] ;
 wire \srfp.register_file[3][16] ;
 wire \srfp.register_file[3][17] ;
 wire \srfp.register_file[3][18] ;
 wire \srfp.register_file[3][19] ;
 wire \srfp.register_file[3][1] ;
 wire \srfp.register_file[3][20] ;
 wire \srfp.register_file[3][21] ;
 wire \srfp.register_file[3][22] ;
 wire \srfp.register_file[3][23] ;
 wire \srfp.register_file[3][24] ;
 wire \srfp.register_file[3][25] ;
 wire \srfp.register_file[3][26] ;
 wire \srfp.register_file[3][27] ;
 wire \srfp.register_file[3][28] ;
 wire \srfp.register_file[3][29] ;
 wire \srfp.register_file[3][2] ;
 wire \srfp.register_file[3][30] ;
 wire \srfp.register_file[3][31] ;
 wire \srfp.register_file[3][3] ;
 wire \srfp.register_file[3][4] ;
 wire \srfp.register_file[3][5] ;
 wire \srfp.register_file[3][6] ;
 wire \srfp.register_file[3][7] ;
 wire \srfp.register_file[3][8] ;
 wire \srfp.register_file[3][9] ;
 wire \srfp.register_file[4][0] ;
 wire \srfp.register_file[4][10] ;
 wire \srfp.register_file[4][11] ;
 wire \srfp.register_file[4][12] ;
 wire \srfp.register_file[4][13] ;
 wire \srfp.register_file[4][14] ;
 wire \srfp.register_file[4][15] ;
 wire \srfp.register_file[4][16] ;
 wire \srfp.register_file[4][17] ;
 wire \srfp.register_file[4][18] ;
 wire \srfp.register_file[4][19] ;
 wire \srfp.register_file[4][1] ;
 wire \srfp.register_file[4][20] ;
 wire \srfp.register_file[4][21] ;
 wire \srfp.register_file[4][22] ;
 wire \srfp.register_file[4][23] ;
 wire \srfp.register_file[4][24] ;
 wire \srfp.register_file[4][25] ;
 wire \srfp.register_file[4][26] ;
 wire \srfp.register_file[4][27] ;
 wire \srfp.register_file[4][28] ;
 wire \srfp.register_file[4][29] ;
 wire \srfp.register_file[4][2] ;
 wire \srfp.register_file[4][30] ;
 wire \srfp.register_file[4][31] ;
 wire \srfp.register_file[4][3] ;
 wire \srfp.register_file[4][4] ;
 wire \srfp.register_file[4][5] ;
 wire \srfp.register_file[4][6] ;
 wire \srfp.register_file[4][7] ;
 wire \srfp.register_file[4][8] ;
 wire \srfp.register_file[4][9] ;
 wire \srfp.register_file[5][0] ;
 wire \srfp.register_file[5][10] ;
 wire \srfp.register_file[5][11] ;
 wire \srfp.register_file[5][12] ;
 wire \srfp.register_file[5][13] ;
 wire \srfp.register_file[5][14] ;
 wire \srfp.register_file[5][15] ;
 wire \srfp.register_file[5][16] ;
 wire \srfp.register_file[5][17] ;
 wire \srfp.register_file[5][18] ;
 wire \srfp.register_file[5][19] ;
 wire \srfp.register_file[5][1] ;
 wire \srfp.register_file[5][20] ;
 wire \srfp.register_file[5][21] ;
 wire \srfp.register_file[5][22] ;
 wire \srfp.register_file[5][23] ;
 wire \srfp.register_file[5][24] ;
 wire \srfp.register_file[5][25] ;
 wire \srfp.register_file[5][26] ;
 wire \srfp.register_file[5][27] ;
 wire \srfp.register_file[5][28] ;
 wire \srfp.register_file[5][29] ;
 wire \srfp.register_file[5][2] ;
 wire \srfp.register_file[5][30] ;
 wire \srfp.register_file[5][31] ;
 wire \srfp.register_file[5][3] ;
 wire \srfp.register_file[5][4] ;
 wire \srfp.register_file[5][5] ;
 wire \srfp.register_file[5][6] ;
 wire \srfp.register_file[5][7] ;
 wire \srfp.register_file[5][8] ;
 wire \srfp.register_file[5][9] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\srfp.register_file[3][16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\srfp.register_file[4][21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0064_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0486_));
 sky130_fd_sc_hd__decap_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__inv_2 _0511_ (.A(net126),
    .Y(_0000_));
 sky130_fd_sc_hd__or4b_2 _0512_ (.A(net6),
    .B(net5),
    .C(net7),
    .D_N(net40),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _0513_ (.A0(net32),
    .A1(\srfp.register_file[0][31] ),
    .S(net120),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _0514_ (.A0(net31),
    .A1(\srfp.register_file[0][30] ),
    .S(net122),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _0515_ (.A0(net29),
    .A1(\srfp.register_file[0][29] ),
    .S(net120),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _0516_ (.A0(net28),
    .A1(\srfp.register_file[0][28] ),
    .S(net120),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _0517_ (.A0(net27),
    .A1(\srfp.register_file[0][27] ),
    .S(net122),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _0518_ (.A0(net26),
    .A1(\srfp.register_file[0][26] ),
    .S(net123),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _0519_ (.A0(net25),
    .A1(\srfp.register_file[0][25] ),
    .S(net122),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _0520_ (.A0(net24),
    .A1(\srfp.register_file[0][24] ),
    .S(net121),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _0521_ (.A0(net23),
    .A1(\srfp.register_file[0][23] ),
    .S(net122),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _0522_ (.A0(net22),
    .A1(\srfp.register_file[0][22] ),
    .S(net120),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _0523_ (.A0(net21),
    .A1(\srfp.register_file[0][21] ),
    .S(net122),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _0524_ (.A0(net20),
    .A1(\srfp.register_file[0][20] ),
    .S(net121),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _0525_ (.A0(net18),
    .A1(\srfp.register_file[0][19] ),
    .S(net120),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _0526_ (.A0(net17),
    .A1(\srfp.register_file[0][18] ),
    .S(net123),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _0527_ (.A0(net16),
    .A1(\srfp.register_file[0][17] ),
    .S(net122),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _0528_ (.A0(net15),
    .A1(\srfp.register_file[0][16] ),
    .S(net121),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _0529_ (.A0(net14),
    .A1(\srfp.register_file[0][15] ),
    .S(net120),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _0530_ (.A0(net13),
    .A1(\srfp.register_file[0][14] ),
    .S(net120),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _0531_ (.A0(net12),
    .A1(\srfp.register_file[0][13] ),
    .S(net121),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _0532_ (.A0(net11),
    .A1(\srfp.register_file[0][12] ),
    .S(net121),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _0533_ (.A0(net10),
    .A1(\srfp.register_file[0][11] ),
    .S(net123),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _0534_ (.A0(net9),
    .A1(\srfp.register_file[0][10] ),
    .S(net121),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _0535_ (.A0(net39),
    .A1(\srfp.register_file[0][9] ),
    .S(net122),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _0536_ (.A0(net38),
    .A1(\srfp.register_file[0][8] ),
    .S(net120),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _0537_ (.A0(net37),
    .A1(\srfp.register_file[0][7] ),
    .S(net120),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _0538_ (.A0(net36),
    .A1(\srfp.register_file[0][6] ),
    .S(net121),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _0539_ (.A0(net35),
    .A1(\srfp.register_file[0][5] ),
    .S(net122),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _0540_ (.A0(net34),
    .A1(\srfp.register_file[0][4] ),
    .S(net122),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _0541_ (.A0(net33),
    .A1(\srfp.register_file[0][3] ),
    .S(net123),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _0542_ (.A0(net30),
    .A1(\srfp.register_file[0][2] ),
    .S(net121),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _0543_ (.A0(net19),
    .A1(\srfp.register_file[0][1] ),
    .S(net122),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _0544_ (.A0(net8),
    .A1(\srfp.register_file[0][0] ),
    .S(net120),
    .X(_0352_));
 sky130_fd_sc_hd__or4bb_1 _0545_ (.A(net6),
    .B(net7),
    .C_N(net40),
    .D_N(net5),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_4 _0546_ (.A0(net32),
    .A1(\srfp.register_file[1][31] ),
    .S(net116),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _0547_ (.A0(net31),
    .A1(\srfp.register_file[1][30] ),
    .S(net118),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _0548_ (.A0(net29),
    .A1(\srfp.register_file[1][29] ),
    .S(net116),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _0549_ (.A0(net28),
    .A1(\srfp.register_file[1][28] ),
    .S(net118),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _0550_ (.A0(net27),
    .A1(\srfp.register_file[1][27] ),
    .S(net116),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _0551_ (.A0(net26),
    .A1(\srfp.register_file[1][26] ),
    .S(net117),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _0552_ (.A0(net25),
    .A1(\srfp.register_file[1][25] ),
    .S(net118),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _0553_ (.A0(net24),
    .A1(\srfp.register_file[1][24] ),
    .S(net117),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _0554_ (.A0(net23),
    .A1(\srfp.register_file[1][23] ),
    .S(net118),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _0555_ (.A0(net22),
    .A1(\srfp.register_file[1][22] ),
    .S(net117),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _0556_ (.A0(net21),
    .A1(\srfp.register_file[1][21] ),
    .S(net118),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _0557_ (.A0(net20),
    .A1(\srfp.register_file[1][20] ),
    .S(net116),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _0558_ (.A0(net18),
    .A1(\srfp.register_file[1][19] ),
    .S(net116),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _0559_ (.A0(net17),
    .A1(\srfp.register_file[1][18] ),
    .S(net118),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _0560_ (.A0(net16),
    .A1(\srfp.register_file[1][17] ),
    .S(net119),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _0561_ (.A0(net15),
    .A1(\srfp.register_file[1][16] ),
    .S(net117),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _0562_ (.A0(net14),
    .A1(\srfp.register_file[1][15] ),
    .S(net118),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _0563_ (.A0(net13),
    .A1(\srfp.register_file[1][14] ),
    .S(net116),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _0564_ (.A0(net12),
    .A1(\srfp.register_file[1][13] ),
    .S(net118),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _0565_ (.A0(net11),
    .A1(\srfp.register_file[1][12] ),
    .S(net117),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _0566_ (.A0(net10),
    .A1(\srfp.register_file[1][11] ),
    .S(net117),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _0567_ (.A0(net9),
    .A1(\srfp.register_file[1][10] ),
    .S(net116),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _0568_ (.A0(net39),
    .A1(\srfp.register_file[1][9] ),
    .S(net119),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_2 _0569_ (.A0(net38),
    .A1(\srfp.register_file[1][8] ),
    .S(net117),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _0570_ (.A0(net37),
    .A1(\srfp.register_file[1][7] ),
    .S(net118),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _0571_ (.A0(net36),
    .A1(\srfp.register_file[1][6] ),
    .S(net116),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _0572_ (.A0(net35),
    .A1(\srfp.register_file[1][5] ),
    .S(net116),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _0573_ (.A0(net34),
    .A1(\srfp.register_file[1][4] ),
    .S(net118),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _0574_ (.A0(net33),
    .A1(\srfp.register_file[1][3] ),
    .S(net119),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_2 _0575_ (.A0(net30),
    .A1(\srfp.register_file[1][2] ),
    .S(net117),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _0576_ (.A0(net19),
    .A1(\srfp.register_file[1][1] ),
    .S(net119),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _0577_ (.A0(net8),
    .A1(\srfp.register_file[1][0] ),
    .S(net116),
    .X(_0320_));
 sky130_fd_sc_hd__or4bb_4 _0578_ (.A(net5),
    .B(net7),
    .C_N(net40),
    .D_N(net6),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _0579_ (.A0(net32),
    .A1(\srfp.register_file[2][31] ),
    .S(net112),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _0580_ (.A0(net31),
    .A1(\srfp.register_file[2][30] ),
    .S(net112),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _0581_ (.A0(net29),
    .A1(\srfp.register_file[2][29] ),
    .S(net115),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _0582_ (.A0(net28),
    .A1(\srfp.register_file[2][28] ),
    .S(net115),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _0583_ (.A0(net27),
    .A1(\srfp.register_file[2][27] ),
    .S(net112),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _0584_ (.A0(net26),
    .A1(\srfp.register_file[2][26] ),
    .S(net115),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _0585_ (.A0(net25),
    .A1(\srfp.register_file[2][25] ),
    .S(net114),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _0586_ (.A0(net24),
    .A1(\srfp.register_file[2][24] ),
    .S(net113),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_2 _0587_ (.A0(net23),
    .A1(\srfp.register_file[2][23] ),
    .S(net115),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _0588_ (.A0(net22),
    .A1(\srfp.register_file[2][22] ),
    .S(net113),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _0589_ (.A0(net21),
    .A1(\srfp.register_file[2][21] ),
    .S(net114),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _0590_ (.A0(net20),
    .A1(\srfp.register_file[2][20] ),
    .S(net114),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _0591_ (.A0(net18),
    .A1(\srfp.register_file[2][19] ),
    .S(net114),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _0592_ (.A0(net17),
    .A1(\srfp.register_file[2][18] ),
    .S(net114),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _0593_ (.A0(net16),
    .A1(\srfp.register_file[2][17] ),
    .S(net115),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _0594_ (.A0(net15),
    .A1(\srfp.register_file[2][16] ),
    .S(net115),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _0595_ (.A0(net14),
    .A1(\srfp.register_file[2][15] ),
    .S(net114),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _0596_ (.A0(net13),
    .A1(\srfp.register_file[2][14] ),
    .S(net112),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _0597_ (.A0(net12),
    .A1(\srfp.register_file[2][13] ),
    .S(net112),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _0598_ (.A0(net11),
    .A1(\srfp.register_file[2][12] ),
    .S(net113),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _0599_ (.A0(net10),
    .A1(\srfp.register_file[2][11] ),
    .S(net112),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_2 _0600_ (.A0(net9),
    .A1(\srfp.register_file[2][10] ),
    .S(net112),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _0601_ (.A0(net39),
    .A1(\srfp.register_file[2][9] ),
    .S(net112),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _0602_ (.A0(net38),
    .A1(\srfp.register_file[2][8] ),
    .S(net113),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _0603_ (.A0(net37),
    .A1(\srfp.register_file[2][7] ),
    .S(net114),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _0604_ (.A0(net36),
    .A1(\srfp.register_file[2][6] ),
    .S(net112),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _0605_ (.A0(net35),
    .A1(\srfp.register_file[2][5] ),
    .S(net114),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _0606_ (.A0(net34),
    .A1(\srfp.register_file[2][4] ),
    .S(net114),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_4 _0607_ (.A0(net33),
    .A1(\srfp.register_file[2][3] ),
    .S(net115),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _0608_ (.A0(net30),
    .A1(\srfp.register_file[2][2] ),
    .S(net113),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _0609_ (.A0(net19),
    .A1(\srfp.register_file[2][1] ),
    .S(net114),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _0610_ (.A0(net8),
    .A1(\srfp.register_file[2][0] ),
    .S(net112),
    .X(_0288_));
 sky130_fd_sc_hd__and4b_4 _0611_ (.A_N(net7),
    .B(net40),
    .C(net6),
    .D(net5),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _0612_ (.A0(\srfp.register_file[3][31] ),
    .A1(net32),
    .S(net108),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _0613_ (.A0(\srfp.register_file[3][30] ),
    .A1(net31),
    .S(net111),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _0614_ (.A0(\srfp.register_file[3][29] ),
    .A1(net29),
    .S(net108),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _0615_ (.A0(\srfp.register_file[3][28] ),
    .A1(net28),
    .S(net110),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _0616_ (.A0(\srfp.register_file[3][27] ),
    .A1(net27),
    .S(net108),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _0617_ (.A0(\srfp.register_file[3][26] ),
    .A1(net26),
    .S(net111),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _0618_ (.A0(\srfp.register_file[3][25] ),
    .A1(net25),
    .S(net110),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _0619_ (.A0(\srfp.register_file[3][24] ),
    .A1(net24),
    .S(net110),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _0620_ (.A0(\srfp.register_file[3][23] ),
    .A1(net23),
    .S(net111),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _0621_ (.A0(\srfp.register_file[3][22] ),
    .A1(net22),
    .S(net109),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _0622_ (.A0(\srfp.register_file[3][21] ),
    .A1(net21),
    .S(net110),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _0623_ (.A0(\srfp.register_file[3][20] ),
    .A1(net20),
    .S(net110),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_2 _0624_ (.A0(\srfp.register_file[3][19] ),
    .A1(net18),
    .S(net108),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _0625_ (.A0(\srfp.register_file[3][18] ),
    .A1(net17),
    .S(net110),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _0626_ (.A0(\srfp.register_file[3][17] ),
    .A1(net16),
    .S(net111),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _0627_ (.A0(\srfp.register_file[3][16] ),
    .A1(net15),
    .S(net110),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _0628_ (.A0(\srfp.register_file[3][15] ),
    .A1(net14),
    .S(net111),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _0629_ (.A0(\srfp.register_file[3][14] ),
    .A1(net13),
    .S(net108),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(\srfp.register_file[3][13] ),
    .A1(net12),
    .S(net108),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _0631_ (.A0(\srfp.register_file[3][12] ),
    .A1(net11),
    .S(net109),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _0632_ (.A0(\srfp.register_file[3][11] ),
    .A1(net10),
    .S(net109),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _0633_ (.A0(\srfp.register_file[3][10] ),
    .A1(net9),
    .S(net110),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _0634_ (.A0(\srfp.register_file[3][9] ),
    .A1(net39),
    .S(net111),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _0635_ (.A0(\srfp.register_file[3][8] ),
    .A1(net38),
    .S(net109),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(\srfp.register_file[3][7] ),
    .A1(net37),
    .S(net108),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_4 _0637_ (.A0(\srfp.register_file[3][6] ),
    .A1(net36),
    .S(net111),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _0638_ (.A0(\srfp.register_file[3][5] ),
    .A1(net35),
    .S(net108),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _0639_ (.A0(\srfp.register_file[3][4] ),
    .A1(net34),
    .S(net110),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _0640_ (.A0(\srfp.register_file[3][3] ),
    .A1(net33),
    .S(net110),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _0641_ (.A0(\srfp.register_file[3][2] ),
    .A1(net30),
    .S(net109),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _0642_ (.A0(\srfp.register_file[3][1] ),
    .A1(net19),
    .S(net108),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_2 _0643_ (.A0(\srfp.register_file[3][0] ),
    .A1(net8),
    .S(net108),
    .X(_0256_));
 sky130_fd_sc_hd__or4bb_2 _0644_ (.A(net6),
    .B(net5),
    .C_N(net7),
    .D_N(net40),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _0645_ (.A0(net32),
    .A1(\srfp.register_file[4][31] ),
    .S(net104),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(net31),
    .A1(\srfp.register_file[4][30] ),
    .S(net105),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _0647_ (.A0(net29),
    .A1(\srfp.register_file[4][29] ),
    .S(net104),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_2 _0648_ (.A0(net28),
    .A1(\srfp.register_file[4][28] ),
    .S(net105),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(net27),
    .A1(\srfp.register_file[4][27] ),
    .S(net105),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0650_ (.A0(net26),
    .A1(\srfp.register_file[4][26] ),
    .S(net106),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_2 _0651_ (.A0(net25),
    .A1(\srfp.register_file[4][25] ),
    .S(net106),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _0652_ (.A0(net24),
    .A1(\srfp.register_file[4][24] ),
    .S(net104),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _0653_ (.A0(net23),
    .A1(\srfp.register_file[4][23] ),
    .S(net106),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _0654_ (.A0(net22),
    .A1(\srfp.register_file[4][22] ),
    .S(net107),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_2 _0655_ (.A0(net21),
    .A1(\srfp.register_file[4][21] ),
    .S(net106),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _0656_ (.A0(net20),
    .A1(\srfp.register_file[4][20] ),
    .S(net104),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _0657_ (.A0(net18),
    .A1(\srfp.register_file[4][19] ),
    .S(net104),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _0658_ (.A0(net17),
    .A1(\srfp.register_file[4][18] ),
    .S(net106),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _0659_ (.A0(net16),
    .A1(\srfp.register_file[4][17] ),
    .S(net105),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _0660_ (.A0(net15),
    .A1(\srfp.register_file[4][16] ),
    .S(net107),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _0661_ (.A0(net14),
    .A1(\srfp.register_file[4][15] ),
    .S(net105),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0662_ (.A0(net13),
    .A1(\srfp.register_file[4][14] ),
    .S(net104),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _0663_ (.A0(net12),
    .A1(\srfp.register_file[4][13] ),
    .S(net104),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0664_ (.A0(net11),
    .A1(\srfp.register_file[4][12] ),
    .S(net104),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _0665_ (.A0(net10),
    .A1(\srfp.register_file[4][11] ),
    .S(net106),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _0666_ (.A0(net9),
    .A1(\srfp.register_file[4][10] ),
    .S(net104),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _0667_ (.A0(net39),
    .A1(\srfp.register_file[4][9] ),
    .S(net106),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_2 _0668_ (.A0(net38),
    .A1(\srfp.register_file[4][8] ),
    .S(net107),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _0669_ (.A0(net37),
    .A1(\srfp.register_file[4][7] ),
    .S(net105),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _0670_ (.A0(net36),
    .A1(\srfp.register_file[4][6] ),
    .S(net106),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _0671_ (.A0(net35),
    .A1(\srfp.register_file[4][5] ),
    .S(net105),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _0672_ (.A0(net34),
    .A1(\srfp.register_file[4][4] ),
    .S(net105),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _0673_ (.A0(net33),
    .A1(\srfp.register_file[4][3] ),
    .S(net105),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _0674_ (.A0(net30),
    .A1(\srfp.register_file[4][2] ),
    .S(net107),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _0675_ (.A0(net19),
    .A1(\srfp.register_file[4][1] ),
    .S(net105),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _0676_ (.A0(net8),
    .A1(\srfp.register_file[4][0] ),
    .S(net104),
    .X(_0224_));
 sky130_fd_sc_hd__and4b_4 _0677_ (.A_N(net6),
    .B(net5),
    .C(net7),
    .D(net40),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _0678_ (.A0(\srfp.register_file[5][31] ),
    .A1(net32),
    .S(net101),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _0679_ (.A0(\srfp.register_file[5][30] ),
    .A1(net31),
    .S(net102),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _0680_ (.A0(\srfp.register_file[5][29] ),
    .A1(net29),
    .S(net100),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _0681_ (.A0(\srfp.register_file[5][28] ),
    .A1(net28),
    .S(net102),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _0682_ (.A0(\srfp.register_file[5][27] ),
    .A1(net27),
    .S(net100),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _0683_ (.A0(\srfp.register_file[5][26] ),
    .A1(net26),
    .S(net103),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _0684_ (.A0(\srfp.register_file[5][25] ),
    .A1(net25),
    .S(net102),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _0685_ (.A0(\srfp.register_file[5][24] ),
    .A1(net24),
    .S(net100),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _0686_ (.A0(\srfp.register_file[5][23] ),
    .A1(net23),
    .S(net102),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(\srfp.register_file[5][22] ),
    .A1(net22),
    .S(net100),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _0688_ (.A0(\srfp.register_file[5][21] ),
    .A1(net21),
    .S(net103),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _0689_ (.A0(\srfp.register_file[5][20] ),
    .A1(net20),
    .S(net100),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _0690_ (.A0(\srfp.register_file[5][19] ),
    .A1(net18),
    .S(net101),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _0691_ (.A0(\srfp.register_file[5][18] ),
    .A1(net17),
    .S(net103),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_2 _0692_ (.A0(\srfp.register_file[5][17] ),
    .A1(net16),
    .S(net103),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _0693_ (.A0(\srfp.register_file[5][16] ),
    .A1(net15),
    .S(net102),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _0694_ (.A0(\srfp.register_file[5][15] ),
    .A1(net14),
    .S(net100),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _0695_ (.A0(\srfp.register_file[5][14] ),
    .A1(net13),
    .S(net100),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _0696_ (.A0(\srfp.register_file[5][13] ),
    .A1(net12),
    .S(net101),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _0697_ (.A0(\srfp.register_file[5][12] ),
    .A1(net11),
    .S(net100),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _0698_ (.A0(\srfp.register_file[5][11] ),
    .A1(net10),
    .S(net103),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _0699_ (.A0(\srfp.register_file[5][10] ),
    .A1(net9),
    .S(net102),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _0700_ (.A0(\srfp.register_file[5][9] ),
    .A1(net39),
    .S(net102),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _0701_ (.A0(\srfp.register_file[5][8] ),
    .A1(net38),
    .S(net100),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _0702_ (.A0(\srfp.register_file[5][7] ),
    .A1(net37),
    .S(net103),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _0703_ (.A0(\srfp.register_file[5][6] ),
    .A1(net36),
    .S(net101),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _0704_ (.A0(\srfp.register_file[5][5] ),
    .A1(net35),
    .S(net102),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _0705_ (.A0(\srfp.register_file[5][4] ),
    .A1(net34),
    .S(net102),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _0706_ (.A0(\srfp.register_file[5][3] ),
    .A1(net33),
    .S(net103),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(\srfp.register_file[5][2] ),
    .A1(net30),
    .S(net101),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _0708_ (.A0(\srfp.register_file[5][1] ),
    .A1(net19),
    .S(net102),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _0709_ (.A0(\srfp.register_file[5][0] ),
    .A1(net8),
    .S(net100),
    .X(_0192_));
 sky130_fd_sc_hd__nor3b_4 _0710_ (.A(net152),
    .B(net150),
    .C_N(net154),
    .Y(_0390_));
 sky130_fd_sc_hd__and2_1 _0711_ (.A(\srfp.register_file[1][0] ),
    .B(net96),
    .X(_0391_));
 sky130_fd_sc_hd__and3b_4 _0712_ (.A_N(net152),
    .B(net154),
    .C(net150),
    .X(_0392_));
 sky130_fd_sc_hd__nand2b_2 _0713_ (.A_N(net150),
    .B(net152),
    .Y(_0393_));
 sky130_fd_sc_hd__nor3b_4 _0714_ (.A(net154),
    .B(net150),
    .C_N(net152),
    .Y(_0394_));
 sky130_fd_sc_hd__a22o_1 _0715_ (.A1(\srfp.register_file[5][0] ),
    .A2(net92),
    .B1(net84),
    .B2(\srfp.register_file[2][0] ),
    .X(_0395_));
 sky130_fd_sc_hd__nor3b_1 _0716_ (.A(net152),
    .B(net154),
    .C_N(net150),
    .Y(_0396_));
 sky130_fd_sc_hd__and3b_2 _0717_ (.A_N(net150),
    .B(net154),
    .C(net152),
    .X(_0397_));
 sky130_fd_sc_hd__o21bai_4 _0718_ (.A1(net154),
    .A2(net150),
    .B1_N(net152),
    .Y(_0398_));
 sky130_fd_sc_hd__and3_1 _0719_ (.A(\srfp.register_file[0][0] ),
    .B(net88),
    .C(net73),
    .X(_0399_));
 sky130_fd_sc_hd__a22o_1 _0720_ (.A1(\srfp.register_file[4][0] ),
    .A2(net81),
    .B1(net77),
    .B2(\srfp.register_file[3][0] ),
    .X(_0400_));
 sky130_fd_sc_hd__or4_1 _0721_ (.A(_0391_),
    .B(_0395_),
    .C(_0399_),
    .D(_0400_),
    .X(net41));
 sky130_fd_sc_hd__and2_1 _0722_ (.A(\srfp.register_file[1][1] ),
    .B(net99),
    .X(_0401_));
 sky130_fd_sc_hd__a22o_1 _0723_ (.A1(\srfp.register_file[5][1] ),
    .A2(net94),
    .B1(net86),
    .B2(\srfp.register_file[2][1] ),
    .X(_0402_));
 sky130_fd_sc_hd__and3_1 _0724_ (.A(\srfp.register_file[0][1] ),
    .B(net90),
    .C(net75),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _0725_ (.A1(\srfp.register_file[4][1] ),
    .A2(net82),
    .B1(net79),
    .B2(\srfp.register_file[3][1] ),
    .X(_0404_));
 sky130_fd_sc_hd__or4_1 _0726_ (.A(_0401_),
    .B(_0402_),
    .C(_0403_),
    .D(_0404_),
    .X(net52));
 sky130_fd_sc_hd__and4bb_1 _0727_ (.A_N(net152),
    .B_N(net154),
    .C(net150),
    .D(\srfp.register_file[4][2] ),
    .X(_0405_));
 sky130_fd_sc_hd__a221o_1 _0728_ (.A1(\srfp.register_file[1][2] ),
    .A2(net97),
    .B1(net85),
    .B2(\srfp.register_file[2][2] ),
    .C1(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__and3_1 _0729_ (.A(\srfp.register_file[0][2] ),
    .B(net89),
    .C(net74),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_1 _0730_ (.A1(\srfp.register_file[5][2] ),
    .A2(net93),
    .B1(net78),
    .B2(\srfp.register_file[3][2] ),
    .X(_0408_));
 sky130_fd_sc_hd__or3_1 _0731_ (.A(_0406_),
    .B(_0407_),
    .C(_0408_),
    .X(net63));
 sky130_fd_sc_hd__a22o_1 _0732_ (.A1(\srfp.register_file[5][3] ),
    .A2(net95),
    .B1(net87),
    .B2(\srfp.register_file[2][3] ),
    .X(_0409_));
 sky130_fd_sc_hd__a22o_1 _0733_ (.A1(\srfp.register_file[1][3] ),
    .A2(net99),
    .B1(net80),
    .B2(\srfp.register_file[3][3] ),
    .X(_0410_));
 sky130_fd_sc_hd__and3_1 _0734_ (.A(\srfp.register_file[0][3] ),
    .B(net91),
    .C(net76),
    .X(_0411_));
 sky130_fd_sc_hd__a2111o_1 _0735_ (.A1(\srfp.register_file[4][3] ),
    .A2(net82),
    .B1(_0409_),
    .C1(_0410_),
    .D1(_0411_),
    .X(net66));
 sky130_fd_sc_hd__and2_1 _0736_ (.A(\srfp.register_file[1][4] ),
    .B(net98),
    .X(_0412_));
 sky130_fd_sc_hd__a22o_1 _0737_ (.A1(\srfp.register_file[5][4] ),
    .A2(net94),
    .B1(net86),
    .B2(\srfp.register_file[2][4] ),
    .X(_0413_));
 sky130_fd_sc_hd__and3_1 _0738_ (.A(\srfp.register_file[0][4] ),
    .B(net90),
    .C(net75),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _0739_ (.A1(\srfp.register_file[4][4] ),
    .A2(net82),
    .B1(net79),
    .B2(\srfp.register_file[3][4] ),
    .X(_0415_));
 sky130_fd_sc_hd__or4_2 _0740_ (.A(_0412_),
    .B(_0413_),
    .C(_0414_),
    .D(_0415_),
    .X(net67));
 sky130_fd_sc_hd__a22o_1 _0741_ (.A1(\srfp.register_file[5][5] ),
    .A2(net94),
    .B1(net87),
    .B2(\srfp.register_file[2][5] ),
    .X(_0416_));
 sky130_fd_sc_hd__a22o_1 _0742_ (.A1(\srfp.register_file[1][5] ),
    .A2(net98),
    .B1(net79),
    .B2(\srfp.register_file[3][5] ),
    .X(_0417_));
 sky130_fd_sc_hd__and3_1 _0743_ (.A(\srfp.register_file[0][5] ),
    .B(net90),
    .C(net75),
    .X(_0418_));
 sky130_fd_sc_hd__a2111o_2 _0744_ (.A1(\srfp.register_file[4][5] ),
    .A2(net82),
    .B1(_0416_),
    .C1(_0417_),
    .D1(_0418_),
    .X(net68));
 sky130_fd_sc_hd__a22o_1 _0745_ (.A1(\srfp.register_file[5][6] ),
    .A2(net92),
    .B1(net84),
    .B2(\srfp.register_file[2][6] ),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _0746_ (.A1(\srfp.register_file[1][6] ),
    .A2(net96),
    .B1(net78),
    .B2(\srfp.register_file[3][6] ),
    .X(_0420_));
 sky130_fd_sc_hd__and3_1 _0747_ (.A(\srfp.register_file[0][6] ),
    .B(net89),
    .C(net74),
    .X(_0421_));
 sky130_fd_sc_hd__a2111o_2 _0748_ (.A1(\srfp.register_file[4][6] ),
    .A2(net81),
    .B1(_0419_),
    .C1(_0420_),
    .D1(_0421_),
    .X(net69));
 sky130_fd_sc_hd__and4bb_1 _0749_ (.A_N(net153),
    .B_N(net154),
    .C(net151),
    .D(\srfp.register_file[4][7] ),
    .X(_0422_));
 sky130_fd_sc_hd__a221o_1 _0750_ (.A1(\srfp.register_file[1][7] ),
    .A2(net98),
    .B1(net86),
    .B2(\srfp.register_file[2][7] ),
    .C1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__and3_1 _0751_ (.A(\srfp.register_file[0][7] ),
    .B(net88),
    .C(net73),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _0752_ (.A1(\srfp.register_file[5][7] ),
    .A2(net92),
    .B1(net77),
    .B2(\srfp.register_file[3][7] ),
    .X(_0425_));
 sky130_fd_sc_hd__or3_1 _0753_ (.A(_0423_),
    .B(_0424_),
    .C(_0425_),
    .X(net70));
 sky130_fd_sc_hd__a22o_1 _0754_ (.A1(\srfp.register_file[5][8] ),
    .A2(net92),
    .B1(net84),
    .B2(\srfp.register_file[2][8] ),
    .X(_0426_));
 sky130_fd_sc_hd__a22o_1 _0755_ (.A1(\srfp.register_file[1][8] ),
    .A2(net96),
    .B1(net77),
    .B2(\srfp.register_file[3][8] ),
    .X(_0427_));
 sky130_fd_sc_hd__and3_1 _0756_ (.A(\srfp.register_file[0][8] ),
    .B(net88),
    .C(net73),
    .X(_0428_));
 sky130_fd_sc_hd__a2111o_1 _0757_ (.A1(\srfp.register_file[4][8] ),
    .A2(net83),
    .B1(_0426_),
    .C1(_0427_),
    .D1(_0428_),
    .X(net71));
 sky130_fd_sc_hd__and2_1 _0758_ (.A(\srfp.register_file[1][9] ),
    .B(net99),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _0759_ (.A1(\srfp.register_file[5][9] ),
    .A2(net95),
    .B1(net87),
    .B2(\srfp.register_file[2][9] ),
    .X(_0430_));
 sky130_fd_sc_hd__and3_1 _0760_ (.A(\srfp.register_file[0][9] ),
    .B(net90),
    .C(net75),
    .X(_0431_));
 sky130_fd_sc_hd__a22o_1 _0761_ (.A1(\srfp.register_file[4][9] ),
    .A2(net83),
    .B1(net80),
    .B2(\srfp.register_file[3][9] ),
    .X(_0432_));
 sky130_fd_sc_hd__or4_4 _0762_ (.A(_0429_),
    .B(_0430_),
    .C(_0431_),
    .D(_0432_),
    .X(net72));
 sky130_fd_sc_hd__a22o_1 _0763_ (.A1(\srfp.register_file[5][10] ),
    .A2(net92),
    .B1(net84),
    .B2(\srfp.register_file[2][10] ),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _0764_ (.A1(\srfp.register_file[1][10] ),
    .A2(net96),
    .B1(net77),
    .B2(\srfp.register_file[3][10] ),
    .X(_0434_));
 sky130_fd_sc_hd__and3_1 _0765_ (.A(\srfp.register_file[0][10] ),
    .B(net88),
    .C(net73),
    .X(_0435_));
 sky130_fd_sc_hd__a2111o_4 _0766_ (.A1(\srfp.register_file[4][10] ),
    .A2(net81),
    .B1(_0433_),
    .C1(_0434_),
    .D1(_0435_),
    .X(net42));
 sky130_fd_sc_hd__a22o_1 _0767_ (.A1(\srfp.register_file[5][11] ),
    .A2(net95),
    .B1(net87),
    .B2(\srfp.register_file[2][11] ),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _0768_ (.A1(\srfp.register_file[1][11] ),
    .A2(net97),
    .B1(net78),
    .B2(\srfp.register_file[3][11] ),
    .X(_0437_));
 sky130_fd_sc_hd__and3_1 _0769_ (.A(\srfp.register_file[0][11] ),
    .B(net91),
    .C(net76),
    .X(_0438_));
 sky130_fd_sc_hd__a2111o_1 _0770_ (.A1(\srfp.register_file[4][11] ),
    .A2(net82),
    .B1(_0436_),
    .C1(_0437_),
    .D1(_0438_),
    .X(net43));
 sky130_fd_sc_hd__a22o_1 _0771_ (.A1(\srfp.register_file[5][12] ),
    .A2(net93),
    .B1(net85),
    .B2(\srfp.register_file[2][12] ),
    .X(_0439_));
 sky130_fd_sc_hd__a22o_1 _0772_ (.A1(\srfp.register_file[1][12] ),
    .A2(net97),
    .B1(net78),
    .B2(\srfp.register_file[3][12] ),
    .X(_0440_));
 sky130_fd_sc_hd__and3_1 _0773_ (.A(\srfp.register_file[0][12] ),
    .B(net88),
    .C(net73),
    .X(_0441_));
 sky130_fd_sc_hd__a2111o_2 _0774_ (.A1(\srfp.register_file[4][12] ),
    .A2(net81),
    .B1(_0439_),
    .C1(_0440_),
    .D1(_0441_),
    .X(net44));
 sky130_fd_sc_hd__a22o_1 _0775_ (.A1(\srfp.register_file[5][13] ),
    .A2(net92),
    .B1(net84),
    .B2(\srfp.register_file[2][13] ),
    .X(_0442_));
 sky130_fd_sc_hd__a22o_1 _0776_ (.A1(\srfp.register_file[1][13] ),
    .A2(net96),
    .B1(net77),
    .B2(\srfp.register_file[3][13] ),
    .X(_0443_));
 sky130_fd_sc_hd__and3_1 _0777_ (.A(\srfp.register_file[0][13] ),
    .B(net88),
    .C(net73),
    .X(_0444_));
 sky130_fd_sc_hd__a2111o_4 _0778_ (.A1(\srfp.register_file[4][13] ),
    .A2(net81),
    .B1(_0442_),
    .C1(_0443_),
    .D1(_0444_),
    .X(net45));
 sky130_fd_sc_hd__and2_1 _0779_ (.A(\srfp.register_file[1][14] ),
    .B(net96),
    .X(_0445_));
 sky130_fd_sc_hd__a22o_1 _0780_ (.A1(\srfp.register_file[5][14] ),
    .A2(net92),
    .B1(net84),
    .B2(\srfp.register_file[2][14] ),
    .X(_0446_));
 sky130_fd_sc_hd__and3_1 _0781_ (.A(\srfp.register_file[0][14] ),
    .B(net88),
    .C(net73),
    .X(_0447_));
 sky130_fd_sc_hd__a22o_1 _0782_ (.A1(\srfp.register_file[4][14] ),
    .A2(net81),
    .B1(net77),
    .B2(\srfp.register_file[3][14] ),
    .X(_0448_));
 sky130_fd_sc_hd__or4_4 _0783_ (.A(_0445_),
    .B(_0446_),
    .C(_0447_),
    .D(_0448_),
    .X(net46));
 sky130_fd_sc_hd__and4bb_1 _0784_ (.A_N(net153),
    .B_N(net1),
    .C(net151),
    .D(\srfp.register_file[4][15] ),
    .X(_0449_));
 sky130_fd_sc_hd__a221o_1 _0785_ (.A1(\srfp.register_file[1][15] ),
    .A2(net98),
    .B1(net86),
    .B2(\srfp.register_file[2][15] ),
    .C1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__and3_1 _0786_ (.A(\srfp.register_file[0][15] ),
    .B(net88),
    .C(net73),
    .X(_0451_));
 sky130_fd_sc_hd__a22o_1 _0787_ (.A1(\srfp.register_file[5][15] ),
    .A2(net94),
    .B1(net79),
    .B2(\srfp.register_file[3][15] ),
    .X(_0452_));
 sky130_fd_sc_hd__or3_2 _0788_ (.A(_0450_),
    .B(_0451_),
    .C(_0452_),
    .X(net47));
 sky130_fd_sc_hd__and2_1 _0789_ (.A(\srfp.register_file[1][16] ),
    .B(net97),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_2 _0790_ (.A1(\srfp.register_file[5][16] ),
    .A2(net95),
    .B1(net87),
    .B2(\srfp.register_file[2][16] ),
    .X(_0454_));
 sky130_fd_sc_hd__and3_1 _0791_ (.A(\srfp.register_file[0][16] ),
    .B(net89),
    .C(net74),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _0792_ (.A1(\srfp.register_file[4][16] ),
    .A2(net81),
    .B1(net78),
    .B2(\srfp.register_file[3][16] ),
    .X(_0456_));
 sky130_fd_sc_hd__or4_2 _0793_ (.A(_0453_),
    .B(_0454_),
    .C(_0455_),
    .D(_0456_),
    .X(net48));
 sky130_fd_sc_hd__and4bb_1 _0794_ (.A_N(net153),
    .B_N(net1),
    .C(net151),
    .D(\srfp.register_file[4][17] ),
    .X(_0457_));
 sky130_fd_sc_hd__a221o_1 _0795_ (.A1(\srfp.register_file[1][17] ),
    .A2(net98),
    .B1(net86),
    .B2(\srfp.register_file[2][17] ),
    .C1(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__and3_1 _0796_ (.A(\srfp.register_file[0][17] ),
    .B(net90),
    .C(net75),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _0797_ (.A1(\srfp.register_file[5][17] ),
    .A2(net95),
    .B1(net80),
    .B2(\srfp.register_file[3][17] ),
    .X(_0460_));
 sky130_fd_sc_hd__or3_1 _0798_ (.A(_0458_),
    .B(_0459_),
    .C(_0460_),
    .X(net49));
 sky130_fd_sc_hd__and4bb_1 _0799_ (.A_N(net153),
    .B_N(net1),
    .C(net151),
    .D(\srfp.register_file[4][18] ),
    .X(_0461_));
 sky130_fd_sc_hd__a221o_1 _0800_ (.A1(\srfp.register_file[1][18] ),
    .A2(net99),
    .B1(net86),
    .B2(\srfp.register_file[2][18] ),
    .C1(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__and3_1 _0801_ (.A(\srfp.register_file[0][18] ),
    .B(net91),
    .C(net76),
    .X(_0463_));
 sky130_fd_sc_hd__a22o_1 _0802_ (.A1(\srfp.register_file[5][18] ),
    .A2(net94),
    .B1(net80),
    .B2(\srfp.register_file[3][18] ),
    .X(_0464_));
 sky130_fd_sc_hd__or3_2 _0803_ (.A(_0462_),
    .B(_0463_),
    .C(_0464_),
    .X(net50));
 sky130_fd_sc_hd__a22o_1 _0804_ (.A1(\srfp.register_file[5][19] ),
    .A2(net93),
    .B1(net85),
    .B2(\srfp.register_file[2][19] ),
    .X(_0465_));
 sky130_fd_sc_hd__a22o_1 _0805_ (.A1(\srfp.register_file[1][19] ),
    .A2(net96),
    .B1(net78),
    .B2(\srfp.register_file[3][19] ),
    .X(_0466_));
 sky130_fd_sc_hd__and3_1 _0806_ (.A(\srfp.register_file[0][19] ),
    .B(net88),
    .C(net73),
    .X(_0467_));
 sky130_fd_sc_hd__a2111o_2 _0807_ (.A1(\srfp.register_file[4][19] ),
    .A2(net83),
    .B1(_0465_),
    .C1(_0466_),
    .D1(_0467_),
    .X(net51));
 sky130_fd_sc_hd__and2_1 _0808_ (.A(\srfp.register_file[1][20] ),
    .B(net98),
    .X(_0468_));
 sky130_fd_sc_hd__a22o_1 _0809_ (.A1(\srfp.register_file[5][20] ),
    .A2(net93),
    .B1(net85),
    .B2(\srfp.register_file[2][20] ),
    .X(_0469_));
 sky130_fd_sc_hd__and3_1 _0810_ (.A(\srfp.register_file[0][20] ),
    .B(net89),
    .C(net74),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _0811_ (.A1(\srfp.register_file[4][20] ),
    .A2(net81),
    .B1(net77),
    .B2(\srfp.register_file[3][20] ),
    .X(_0471_));
 sky130_fd_sc_hd__or4_4 _0812_ (.A(_0468_),
    .B(_0469_),
    .C(_0470_),
    .D(_0471_),
    .X(net53));
 sky130_fd_sc_hd__a22o_1 _0813_ (.A1(\srfp.register_file[5][21] ),
    .A2(net94),
    .B1(net86),
    .B2(\srfp.register_file[2][21] ),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _0814_ (.A1(\srfp.register_file[1][21] ),
    .A2(net99),
    .B1(net80),
    .B2(\srfp.register_file[3][21] ),
    .X(_0473_));
 sky130_fd_sc_hd__and3_1 _0815_ (.A(\srfp.register_file[0][21] ),
    .B(net90),
    .C(net75),
    .X(_0474_));
 sky130_fd_sc_hd__a2111o_2 _0816_ (.A1(\srfp.register_file[4][21] ),
    .A2(net82),
    .B1(_0472_),
    .C1(_0473_),
    .D1(_0474_),
    .X(net54));
 sky130_fd_sc_hd__and4bb_1 _0817_ (.A_N(net152),
    .B_N(net154),
    .C(net150),
    .D(\srfp.register_file[4][22] ),
    .X(_0475_));
 sky130_fd_sc_hd__a221o_1 _0818_ (.A1(\srfp.register_file[1][22] ),
    .A2(net96),
    .B1(net84),
    .B2(\srfp.register_file[2][22] ),
    .C1(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__and3_1 _0819_ (.A(\srfp.register_file[0][22] ),
    .B(net88),
    .C(net73),
    .X(_0477_));
 sky130_fd_sc_hd__a22o_1 _0820_ (.A1(\srfp.register_file[5][22] ),
    .A2(net92),
    .B1(net77),
    .B2(\srfp.register_file[3][22] ),
    .X(_0478_));
 sky130_fd_sc_hd__or3_2 _0821_ (.A(_0476_),
    .B(_0477_),
    .C(_0478_),
    .X(net55));
 sky130_fd_sc_hd__and4bb_1 _0822_ (.A_N(net153),
    .B_N(net1),
    .C(net151),
    .D(\srfp.register_file[4][23] ),
    .X(_0479_));
 sky130_fd_sc_hd__a221o_1 _0823_ (.A1(\srfp.register_file[1][23] ),
    .A2(net99),
    .B1(net87),
    .B2(\srfp.register_file[2][23] ),
    .C1(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__and3_1 _0824_ (.A(\srfp.register_file[0][23] ),
    .B(net91),
    .C(net76),
    .X(_0481_));
 sky130_fd_sc_hd__a22o_1 _0825_ (.A1(\srfp.register_file[5][23] ),
    .A2(net94),
    .B1(net79),
    .B2(\srfp.register_file[3][23] ),
    .X(_0482_));
 sky130_fd_sc_hd__or3_1 _0826_ (.A(_0480_),
    .B(_0481_),
    .C(_0482_),
    .X(net56));
 sky130_fd_sc_hd__and2_1 _0827_ (.A(\srfp.register_file[1][24] ),
    .B(net97),
    .X(_0483_));
 sky130_fd_sc_hd__a22o_1 _0828_ (.A1(\srfp.register_file[5][24] ),
    .A2(net93),
    .B1(net85),
    .B2(\srfp.register_file[2][24] ),
    .X(_0484_));
 sky130_fd_sc_hd__and3_1 _0829_ (.A(\srfp.register_file[0][24] ),
    .B(net89),
    .C(net74),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_2 _0830_ (.A1(\srfp.register_file[4][24] ),
    .A2(net81),
    .B1(net77),
    .B2(\srfp.register_file[3][24] ),
    .X(_0486_));
 sky130_fd_sc_hd__or4_1 _0831_ (.A(_0483_),
    .B(_0484_),
    .C(_0485_),
    .D(_0486_),
    .X(net57));
 sky130_fd_sc_hd__a22o_1 _0832_ (.A1(\srfp.register_file[5][25] ),
    .A2(net94),
    .B1(net86),
    .B2(\srfp.register_file[2][25] ),
    .X(_0487_));
 sky130_fd_sc_hd__a22o_1 _0833_ (.A1(\srfp.register_file[1][25] ),
    .A2(net98),
    .B1(net79),
    .B2(\srfp.register_file[3][25] ),
    .X(_0488_));
 sky130_fd_sc_hd__and3_1 _0834_ (.A(\srfp.register_file[0][25] ),
    .B(net90),
    .C(net75),
    .X(_0489_));
 sky130_fd_sc_hd__a2111o_1 _0835_ (.A1(\srfp.register_file[4][25] ),
    .A2(net82),
    .B1(_0487_),
    .C1(_0488_),
    .D1(_0489_),
    .X(net58));
 sky130_fd_sc_hd__a22o_1 _0836_ (.A1(\srfp.register_file[5][26] ),
    .A2(net95),
    .B1(net87),
    .B2(\srfp.register_file[2][26] ),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _0837_ (.A1(\srfp.register_file[1][26] ),
    .A2(net98),
    .B1(net79),
    .B2(\srfp.register_file[3][26] ),
    .X(_0491_));
 sky130_fd_sc_hd__and3_1 _0838_ (.A(\srfp.register_file[0][26] ),
    .B(net91),
    .C(net76),
    .X(_0492_));
 sky130_fd_sc_hd__a2111o_2 _0839_ (.A1(\srfp.register_file[4][26] ),
    .A2(net83),
    .B1(_0490_),
    .C1(_0491_),
    .D1(_0492_),
    .X(net59));
 sky130_fd_sc_hd__a22o_1 _0840_ (.A1(\srfp.register_file[5][27] ),
    .A2(net92),
    .B1(net84),
    .B2(\srfp.register_file[2][27] ),
    .X(_0493_));
 sky130_fd_sc_hd__a22o_1 _0841_ (.A1(\srfp.register_file[1][27] ),
    .A2(net98),
    .B1(net79),
    .B2(\srfp.register_file[3][27] ),
    .X(_0494_));
 sky130_fd_sc_hd__and3_1 _0842_ (.A(\srfp.register_file[0][27] ),
    .B(net90),
    .C(net75),
    .X(_0495_));
 sky130_fd_sc_hd__a2111o_1 _0843_ (.A1(\srfp.register_file[4][27] ),
    .A2(net82),
    .B1(_0493_),
    .C1(_0494_),
    .D1(_0495_),
    .X(net60));
 sky130_fd_sc_hd__and2_1 _0844_ (.A(\srfp.register_file[1][28] ),
    .B(net99),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _0845_ (.A1(\srfp.register_file[5][28] ),
    .A2(net94),
    .B1(net86),
    .B2(\srfp.register_file[2][28] ),
    .X(_0497_));
 sky130_fd_sc_hd__and3_1 _0846_ (.A(\srfp.register_file[0][28] ),
    .B(net90),
    .C(net75),
    .X(_0498_));
 sky130_fd_sc_hd__a22o_1 _0847_ (.A1(\srfp.register_file[4][28] ),
    .A2(net82),
    .B1(net79),
    .B2(\srfp.register_file[3][28] ),
    .X(_0499_));
 sky130_fd_sc_hd__or4_1 _0848_ (.A(_0496_),
    .B(_0497_),
    .C(_0498_),
    .D(_0499_),
    .X(net61));
 sky130_fd_sc_hd__a22o_1 _0849_ (.A1(\srfp.register_file[5][29] ),
    .A2(net92),
    .B1(net84),
    .B2(\srfp.register_file[2][29] ),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _0850_ (.A1(\srfp.register_file[1][29] ),
    .A2(net96),
    .B1(net77),
    .B2(\srfp.register_file[3][29] ),
    .X(_0501_));
 sky130_fd_sc_hd__and3_1 _0851_ (.A(\srfp.register_file[0][29] ),
    .B(net89),
    .C(net74),
    .X(_0502_));
 sky130_fd_sc_hd__a2111o_1 _0852_ (.A1(\srfp.register_file[4][29] ),
    .A2(net81),
    .B1(_0500_),
    .C1(_0501_),
    .D1(_0502_),
    .X(net62));
 sky130_fd_sc_hd__and2_1 _0853_ (.A(\srfp.register_file[1][30] ),
    .B(net98),
    .X(_0503_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(\srfp.register_file[5][30] ),
    .A2(net94),
    .B1(net86),
    .B2(\srfp.register_file[2][30] ),
    .X(_0504_));
 sky130_fd_sc_hd__and3_1 _0855_ (.A(\srfp.register_file[0][30] ),
    .B(net90),
    .C(net75),
    .X(_0505_));
 sky130_fd_sc_hd__a22o_1 _0856_ (.A1(\srfp.register_file[4][30] ),
    .A2(net82),
    .B1(net79),
    .B2(\srfp.register_file[3][30] ),
    .X(_0506_));
 sky130_fd_sc_hd__or4_4 _0857_ (.A(_0503_),
    .B(_0504_),
    .C(_0505_),
    .D(_0506_),
    .X(net64));
 sky130_fd_sc_hd__and4bb_1 _0858_ (.A_N(net152),
    .B_N(net154),
    .C(net150),
    .D(\srfp.register_file[4][31] ),
    .X(_0507_));
 sky130_fd_sc_hd__a221o_1 _0859_ (.A1(\srfp.register_file[1][31] ),
    .A2(net96),
    .B1(net84),
    .B2(\srfp.register_file[2][31] ),
    .C1(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__and3_1 _0860_ (.A(\srfp.register_file[0][31] ),
    .B(net89),
    .C(net74),
    .X(_0509_));
 sky130_fd_sc_hd__a22o_1 _0861_ (.A1(\srfp.register_file[5][31] ),
    .A2(net93),
    .B1(net78),
    .B2(\srfp.register_file[3][31] ),
    .X(_0510_));
 sky130_fd_sc_hd__or3_2 _0862_ (.A(_0508_),
    .B(_0509_),
    .C(_0510_),
    .X(net65));
 sky130_fd_sc_hd__inv_2 _0863_ (.A(net136),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0864_ (.A(net133),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0865_ (.A(net131),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0866_ (.A(net140),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0867_ (.A(net127),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0868_ (.A(net131),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0869_ (.A(net136),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0870_ (.A(net126),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0871_ (.A(net146),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _0872_ (.A(net137),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0873_ (.A(net147),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0874_ (.A(net133),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0875_ (.A(net134),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0876_ (.A(net137),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0877_ (.A(net128),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _0878_ (.A(net144),
    .Y(_0016_));
 sky130_fd_sc_hd__clkinv_2 _0879_ (.A(net146),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _0880_ (.A(net147),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _0881_ (.A(net132),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _0882_ (.A(net134),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _0883_ (.A(net147),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0884_ (.A(net125),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _0885_ (.A(net136),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _0886_ (.A(net131),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0887_ (.A(net127),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _0888_ (.A(net147),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _0889_ (.A(net128),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _0890_ (.A(net140),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0891_ (.A(net126),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _0892_ (.A(net128),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0893_ (.A(net132),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _0894_ (.A(net124),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _0895_ (.A(net141),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _0896_ (.A(net146),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _0897_ (.A(net142),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _0898_ (.A(net140),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _0899_ (.A(net140),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _0900_ (.A(net147),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _0901_ (.A(net138),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _0902_ (.A(net142),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _0903_ (.A(net147),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _0904_ (.A(net127),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _0905_ (.A(net139),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _0906_ (.A(net127),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _0907_ (.A(net126),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _0908_ (.A(net124),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _0909_ (.A(net141),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _0910_ (.A(net133),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _0911_ (.A(net136),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _0912_ (.A(net147),
    .Y(_0050_));
 sky130_fd_sc_hd__clkinv_2 _0913_ (.A(net146),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _0914_ (.A(net134),
    .Y(_0052_));
 sky130_fd_sc_hd__clkinv_2 _0915_ (.A(net147),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _0916_ (.A(net146),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _0917_ (.A(net148),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _0918_ (.A(net128),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _0919_ (.A(net131),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _0920_ (.A(net146),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _0921_ (.A(net141),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _0922_ (.A(net138),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _0923_ (.A(net140),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _0924_ (.A(net136),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _0925_ (.A(net126),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _0926_ (.A(net127),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _0927_ (.A(net124),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _0928_ (.A(net134),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _0929_ (.A(net142),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _0930_ (.A(net140),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _0931_ (.A(net128),
    .Y(_0069_));
 sky130_fd_sc_hd__clkinv_2 _0932_ (.A(net148),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _0933_ (.A(net124),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _0934_ (.A(net133),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _0935_ (.A(net148),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _0936_ (.A(net141),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _0937_ (.A(net134),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _0938_ (.A(net129),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _0939_ (.A(net125),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _0940_ (.A(net126),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _0941_ (.A(net142),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _0942_ (.A(net138),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _0943_ (.A(net146),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _0944_ (.A(net142),
    .Y(_0082_));
 sky130_fd_sc_hd__clkinv_2 _0945_ (.A(net125),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _0946_ (.A(net136),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _0947_ (.A(net142),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _0948_ (.A(net129),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _0949_ (.A(net147),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _0950_ (.A(net137),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _0951_ (.A(net136),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _0952_ (.A(net142),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _0953_ (.A(net138),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _0954_ (.A(net143),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _0955_ (.A(net129),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _0956_ (.A(net146),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _0957_ (.A(net131),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _0958_ (.A(net125),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _0959_ (.A(net137),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _0960_ (.A(net126),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _0961_ (.A(net134),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _0962_ (.A(net137),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _0963_ (.A(net143),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _0964_ (.A(net129),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _0965_ (.A(net140),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _0966_ (.A(net144),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _0967_ (.A(net134),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _0968_ (.A(net140),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _0969_ (.A(net128),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(net133),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _0971_ (.A(net124),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _0972_ (.A(net127),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _0973_ (.A(net142),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _0974_ (.A(net148),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _0975_ (.A(net141),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _0976_ (.A(net139),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _0977_ (.A(net138),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _0978_ (.A(net146),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _0979_ (.A(net138),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _0980_ (.A(net129),
    .Y(_0118_));
 sky130_fd_sc_hd__clkinv_2 _0981_ (.A(net134),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _0982_ (.A(net124),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _0983_ (.A(net124),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _0984_ (.A(net146),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _0985_ (.A(net128),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _0986_ (.A(net137),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _0987_ (.A(net148),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _0988_ (.A(net139),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _0989_ (.A(net124),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(net126),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(net148),
    .Y(_0129_));
 sky130_fd_sc_hd__clkinv_2 _0992_ (.A(net133),
    .Y(_0130_));
 sky130_fd_sc_hd__clkinv_2 _0993_ (.A(net148),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _0994_ (.A(net128),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _0995_ (.A(net131),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _0996_ (.A(net133),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _0997_ (.A(net136),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _0998_ (.A(net129),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _0999_ (.A(net149),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _1000_ (.A(net124),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1001_ (.A(net127),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _1002_ (.A(net133),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _1003_ (.A(net129),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _1004_ (.A(net127),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _1005_ (.A(net138),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1006_ (.A(net131),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _1007_ (.A(net143),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(net136),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1009_ (.A(net125),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _1010_ (.A(net129),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1011_ (.A(net144),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _1012_ (.A(net126),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _1013_ (.A(net142),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _1014_ (.A(net132),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _1015_ (.A(net141),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _1016_ (.A(net127),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _1017_ (.A(net130),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _1018_ (.A(net144),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _1019_ (.A(net125),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _1020_ (.A(net138),
    .Y(_0158_));
 sky130_fd_sc_hd__clkinv_2 _1021_ (.A(net125),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _1022_ (.A(net125),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _1023_ (.A(net140),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _1024_ (.A(net132),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _1025_ (.A(net134),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _1026_ (.A(net137),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _1027_ (.A(net142),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(net131),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _1029_ (.A(net130),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _1030_ (.A(net127),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _1031_ (.A(net148),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _1032_ (.A(net128),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _1033_ (.A(net148),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _1034_ (.A(net133),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _1035_ (.A(net136),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(net124),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _1037_ (.A(net125),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _1038_ (.A(net132),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _1039_ (.A(net143),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _1040_ (.A(net143),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _1041_ (.A(net130),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _1042_ (.A(net131),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _1043_ (.A(net139),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _1044_ (.A(net130),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _1045_ (.A(net149),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _1046_ (.A(net133),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _1047_ (.A(net131),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _1048_ (.A(net149),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(net140),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(net138),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(net130),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(net147),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(net138),
    .Y(_0191_));
 sky130_fd_sc_hd__dfrtp_1 _1054_ (.CLK(clknet_4_4_0_clk),
    .D(_0192_),
    .RESET_B(_0000_),
    .Q(\srfp.register_file[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1055_ (.CLK(clknet_4_8_0_clk),
    .D(_0193_),
    .RESET_B(_0001_),
    .Q(\srfp.register_file[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1056_ (.CLK(clknet_4_7_0_clk),
    .D(_0194_),
    .RESET_B(_0002_),
    .Q(\srfp.register_file[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1057_ (.CLK(clknet_4_13_0_clk),
    .D(_0195_),
    .RESET_B(_0003_),
    .Q(\srfp.register_file[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1058_ (.CLK(clknet_4_10_0_clk),
    .D(_0196_),
    .RESET_B(_0004_),
    .Q(\srfp.register_file[5][4] ));
 sky130_fd_sc_hd__dfrtp_2 _1059_ (.CLK(clknet_4_0_0_clk),
    .D(_0197_),
    .RESET_B(_0005_),
    .Q(\srfp.register_file[5][5] ));
 sky130_fd_sc_hd__dfrtp_2 _1060_ (.CLK(clknet_4_5_0_clk),
    .D(_0198_),
    .RESET_B(_0006_),
    .Q(\srfp.register_file[5][6] ));
 sky130_fd_sc_hd__dfrtp_4 _1061_ (.CLK(clknet_4_9_0_clk),
    .D(_0199_),
    .RESET_B(_0007_),
    .Q(\srfp.register_file[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1062_ (.CLK(clknet_4_1_0_clk),
    .D(_0200_),
    .RESET_B(_0008_),
    .Q(\srfp.register_file[5][8] ));
 sky130_fd_sc_hd__dfrtp_1 _1063_ (.CLK(clknet_4_12_0_clk),
    .D(_0201_),
    .RESET_B(_0009_),
    .Q(\srfp.register_file[5][9] ));
 sky130_fd_sc_hd__dfrtp_1 _1064_ (.CLK(clknet_4_2_0_clk),
    .D(_0202_),
    .RESET_B(_0010_),
    .Q(\srfp.register_file[5][10] ));
 sky130_fd_sc_hd__dfrtp_4 _1065_ (.CLK(clknet_4_15_0_clk),
    .D(_0203_),
    .RESET_B(_0011_),
    .Q(\srfp.register_file[5][11] ));
 sky130_fd_sc_hd__dfrtp_1 _1066_ (.CLK(clknet_4_7_0_clk),
    .D(_0204_),
    .RESET_B(_0012_),
    .Q(\srfp.register_file[5][12] ));
 sky130_fd_sc_hd__dfrtp_2 _1067_ (.CLK(clknet_4_7_0_clk),
    .D(_0205_),
    .RESET_B(_0013_),
    .Q(\srfp.register_file[5][13] ));
 sky130_fd_sc_hd__dfrtp_1 _1068_ (.CLK(clknet_4_0_0_clk),
    .D(_0206_),
    .RESET_B(_0014_),
    .Q(\srfp.register_file[5][14] ));
 sky130_fd_sc_hd__dfrtp_2 _1069_ (.CLK(clknet_4_1_0_clk),
    .D(_0207_),
    .RESET_B(_0015_),
    .Q(\srfp.register_file[5][15] ));
 sky130_fd_sc_hd__dfrtp_1 _1070_ (.CLK(clknet_4_9_0_clk),
    .D(_0208_),
    .RESET_B(_0016_),
    .Q(\srfp.register_file[5][16] ));
 sky130_fd_sc_hd__dfrtp_2 _1071_ (.CLK(clknet_4_2_0_clk),
    .D(_0209_),
    .RESET_B(_0017_),
    .Q(\srfp.register_file[5][17] ));
 sky130_fd_sc_hd__dfrtp_1 _1072_ (.CLK(clknet_4_14_0_clk),
    .D(_0210_),
    .RESET_B(_0018_),
    .Q(\srfp.register_file[5][18] ));
 sky130_fd_sc_hd__dfrtp_2 _1073_ (.CLK(clknet_4_5_0_clk),
    .D(_0211_),
    .RESET_B(_0019_),
    .Q(\srfp.register_file[5][19] ));
 sky130_fd_sc_hd__dfrtp_4 _1074_ (.CLK(clknet_4_7_0_clk),
    .D(_0212_),
    .RESET_B(_0020_),
    .Q(\srfp.register_file[5][20] ));
 sky130_fd_sc_hd__dfrtp_1 _1075_ (.CLK(clknet_4_12_0_clk),
    .D(_0213_),
    .RESET_B(_0021_),
    .Q(\srfp.register_file[5][21] ));
 sky130_fd_sc_hd__dfrtp_1 _1076_ (.CLK(clknet_4_0_0_clk),
    .D(_0214_),
    .RESET_B(_0022_),
    .Q(\srfp.register_file[5][22] ));
 sky130_fd_sc_hd__dfrtp_4 _1077_ (.CLK(clknet_4_8_0_clk),
    .D(_0215_),
    .RESET_B(_0023_),
    .Q(\srfp.register_file[5][23] ));
 sky130_fd_sc_hd__dfrtp_2 _1078_ (.CLK(clknet_4_0_0_clk),
    .D(_0216_),
    .RESET_B(_0024_),
    .Q(\srfp.register_file[5][24] ));
 sky130_fd_sc_hd__dfrtp_1 _1079_ (.CLK(clknet_4_8_0_clk),
    .D(_0217_),
    .RESET_B(_0025_),
    .Q(\srfp.register_file[5][25] ));
 sky130_fd_sc_hd__dfrtp_1 _1080_ (.CLK(clknet_4_15_0_clk),
    .D(_0218_),
    .RESET_B(_0026_),
    .Q(\srfp.register_file[5][26] ));
 sky130_fd_sc_hd__dfrtp_1 _1081_ (.CLK(clknet_4_8_0_clk),
    .D(_0219_),
    .RESET_B(_0027_),
    .Q(\srfp.register_file[5][27] ));
 sky130_fd_sc_hd__dfrtp_1 _1082_ (.CLK(clknet_4_10_0_clk),
    .D(_0220_),
    .RESET_B(_0028_),
    .Q(\srfp.register_file[5][28] ));
 sky130_fd_sc_hd__dfrtp_1 _1083_ (.CLK(clknet_4_0_0_clk),
    .D(_0221_),
    .RESET_B(_0029_),
    .Q(\srfp.register_file[5][29] ));
 sky130_fd_sc_hd__dfrtp_1 _1084_ (.CLK(clknet_4_2_0_clk),
    .D(_0222_),
    .RESET_B(_0030_),
    .Q(\srfp.register_file[5][30] ));
 sky130_fd_sc_hd__dfrtp_1 _1085_ (.CLK(clknet_4_5_0_clk),
    .D(_0223_),
    .RESET_B(_0031_),
    .Q(\srfp.register_file[5][31] ));
 sky130_fd_sc_hd__dfrtp_4 _1086_ (.CLK(clknet_4_2_0_clk),
    .D(_0224_),
    .RESET_B(_0032_),
    .Q(\srfp.register_file[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1087_ (.CLK(clknet_4_10_0_clk),
    .D(_0225_),
    .RESET_B(_0033_),
    .Q(\srfp.register_file[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1088_ (.CLK(clknet_4_5_0_clk),
    .D(_0226_),
    .RESET_B(_0034_),
    .Q(\srfp.register_file[4][2] ));
 sky130_fd_sc_hd__dfrtp_4 _1089_ (.CLK(clknet_4_11_0_clk),
    .D(_0227_),
    .RESET_B(_0035_),
    .Q(\srfp.register_file[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1090_ (.CLK(clknet_4_8_0_clk),
    .D(_0228_),
    .RESET_B(_0036_),
    .Q(\srfp.register_file[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1091_ (.CLK(clknet_4_8_0_clk),
    .D(_0229_),
    .RESET_B(_0037_),
    .Q(\srfp.register_file[4][5] ));
 sky130_fd_sc_hd__dfrtp_2 _1092_ (.CLK(clknet_4_13_0_clk),
    .D(_0230_),
    .RESET_B(_0038_),
    .Q(\srfp.register_file[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1093_ (.CLK(clknet_4_9_0_clk),
    .D(_0231_),
    .RESET_B(_0039_),
    .Q(\srfp.register_file[4][7] ));
 sky130_fd_sc_hd__dfrtp_2 _1094_ (.CLK(clknet_4_12_0_clk),
    .D(_0232_),
    .RESET_B(_0040_),
    .Q(\srfp.register_file[4][8] ));
 sky130_fd_sc_hd__dfrtp_1 _1095_ (.CLK(clknet_4_12_0_clk),
    .D(_0233_),
    .RESET_B(_0041_),
    .Q(\srfp.register_file[4][9] ));
 sky130_fd_sc_hd__dfrtp_1 _1096_ (.CLK(clknet_4_2_0_clk),
    .D(_0234_),
    .RESET_B(_0042_),
    .Q(\srfp.register_file[4][10] ));
 sky130_fd_sc_hd__dfrtp_1 _1097_ (.CLK(clknet_4_13_0_clk),
    .D(_0235_),
    .RESET_B(_0043_),
    .Q(\srfp.register_file[4][11] ));
 sky130_fd_sc_hd__dfrtp_1 _1098_ (.CLK(clknet_4_3_0_clk),
    .D(_0236_),
    .RESET_B(_0044_),
    .Q(\srfp.register_file[4][12] ));
 sky130_fd_sc_hd__dfrtp_1 _1099_ (.CLK(clknet_4_1_0_clk),
    .D(_0237_),
    .RESET_B(_0045_),
    .Q(\srfp.register_file[4][13] ));
 sky130_fd_sc_hd__dfrtp_1 _1100_ (.CLK(clknet_4_0_0_clk),
    .D(_0238_),
    .RESET_B(_0046_),
    .Q(\srfp.register_file[4][14] ));
 sky130_fd_sc_hd__dfrtp_1 _1101_ (.CLK(clknet_4_11_0_clk),
    .D(_0239_),
    .RESET_B(_0047_),
    .Q(\srfp.register_file[4][15] ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_4_7_0_clk),
    .D(_0240_),
    .RESET_B(_0048_),
    .Q(\srfp.register_file[4][16] ));
 sky130_fd_sc_hd__dfrtp_1 _1103_ (.CLK(clknet_4_11_0_clk),
    .D(_0241_),
    .RESET_B(_0049_),
    .Q(\srfp.register_file[4][17] ));
 sky130_fd_sc_hd__dfrtp_4 _1104_ (.CLK(clknet_4_14_0_clk),
    .D(_0242_),
    .RESET_B(_0050_),
    .Q(\srfp.register_file[4][18] ));
 sky130_fd_sc_hd__dfrtp_2 _1105_ (.CLK(clknet_4_0_0_clk),
    .D(_0243_),
    .RESET_B(_0051_),
    .Q(\srfp.register_file[4][19] ));
 sky130_fd_sc_hd__dfrtp_1 _1106_ (.CLK(clknet_4_2_0_clk),
    .D(_0244_),
    .RESET_B(_0052_),
    .Q(\srfp.register_file[4][20] ));
 sky130_fd_sc_hd__dfrtp_2 _1107_ (.CLK(clknet_4_4_0_clk),
    .D(_0245_),
    .RESET_B(_0053_),
    .Q(\srfp.register_file[4][21] ));
 sky130_fd_sc_hd__dfrtp_1 _1108_ (.CLK(clknet_4_7_0_clk),
    .D(_0246_),
    .RESET_B(_0054_),
    .Q(\srfp.register_file[4][22] ));
 sky130_fd_sc_hd__dfrtp_1 _1109_ (.CLK(clknet_4_14_0_clk),
    .D(_0247_),
    .RESET_B(_0055_),
    .Q(\srfp.register_file[4][23] ));
 sky130_fd_sc_hd__dfrtp_1 _1110_ (.CLK(clknet_4_2_0_clk),
    .D(_0248_),
    .RESET_B(_0056_),
    .Q(\srfp.register_file[4][24] ));
 sky130_fd_sc_hd__dfrtp_2 _1111_ (.CLK(clknet_4_10_0_clk),
    .D(_0249_),
    .RESET_B(_0057_),
    .Q(\srfp.register_file[4][25] ));
 sky130_fd_sc_hd__dfrtp_1 _1112_ (.CLK(clknet_4_13_0_clk),
    .D(_0250_),
    .RESET_B(_0058_),
    .Q(\srfp.register_file[4][26] ));
 sky130_fd_sc_hd__dfrtp_4 _1113_ (.CLK(clknet_4_10_0_clk),
    .D(_0251_),
    .RESET_B(_0059_),
    .Q(\srfp.register_file[4][27] ));
 sky130_fd_sc_hd__dfrtp_2 _1114_ (.CLK(clknet_4_1_0_clk),
    .D(_0252_),
    .RESET_B(_0060_),
    .Q(\srfp.register_file[4][28] ));
 sky130_fd_sc_hd__dfrtp_1 _1115_ (.CLK(clknet_4_2_0_clk),
    .D(_0253_),
    .RESET_B(_0061_),
    .Q(\srfp.register_file[4][29] ));
 sky130_fd_sc_hd__dfrtp_1 _1116_ (.CLK(clknet_4_12_0_clk),
    .D(_0254_),
    .RESET_B(_0062_),
    .Q(\srfp.register_file[4][30] ));
 sky130_fd_sc_hd__dfrtp_1 _1117_ (.CLK(clknet_4_4_0_clk),
    .D(_0255_),
    .RESET_B(_0063_),
    .Q(\srfp.register_file[4][31] ));
 sky130_fd_sc_hd__dfrtp_2 _1118_ (.CLK(clknet_4_10_0_clk),
    .D(_0256_),
    .RESET_B(_0064_),
    .Q(\srfp.register_file[3][0] ));
 sky130_fd_sc_hd__dfrtp_4 _1119_ (.CLK(clknet_4_2_0_clk),
    .D(_0257_),
    .RESET_B(_0065_),
    .Q(\srfp.register_file[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_4_7_0_clk),
    .D(_0258_),
    .RESET_B(_0066_),
    .Q(\srfp.register_file[3][2] ));
 sky130_fd_sc_hd__dfrtp_4 _1121_ (.CLK(clknet_4_9_0_clk),
    .D(_0259_),
    .RESET_B(_0067_),
    .Q(\srfp.register_file[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1122_ (.CLK(clknet_4_10_0_clk),
    .D(_0260_),
    .RESET_B(_0068_),
    .Q(\srfp.register_file[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1123_ (.CLK(clknet_4_3_0_clk),
    .D(_0261_),
    .RESET_B(_0069_),
    .Q(\srfp.register_file[3][5] ));
 sky130_fd_sc_hd__dfrtp_2 _1124_ (.CLK(clknet_4_2_0_clk),
    .D(_0262_),
    .RESET_B(_0070_),
    .Q(\srfp.register_file[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1125_ (.CLK(clknet_4_2_0_clk),
    .D(_0263_),
    .RESET_B(_0071_),
    .Q(\srfp.register_file[3][7] ));
 sky130_fd_sc_hd__dfrtp_4 _1126_ (.CLK(clknet_4_7_0_clk),
    .D(_0264_),
    .RESET_B(_0072_),
    .Q(\srfp.register_file[3][8] ));
 sky130_fd_sc_hd__dfrtp_2 _1127_ (.CLK(clknet_4_15_0_clk),
    .D(_0265_),
    .RESET_B(_0073_),
    .Q(\srfp.register_file[3][9] ));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(clknet_4_8_0_clk),
    .D(_0266_),
    .RESET_B(_0074_),
    .Q(\srfp.register_file[3][10] ));
 sky130_fd_sc_hd__dfrtp_1 _1129_ (.CLK(clknet_4_6_0_clk),
    .D(_0267_),
    .RESET_B(_0075_),
    .Q(\srfp.register_file[3][11] ));
 sky130_fd_sc_hd__dfrtp_1 _1130_ (.CLK(clknet_4_6_0_clk),
    .D(_0268_),
    .RESET_B(_0076_),
    .Q(\srfp.register_file[3][12] ));
 sky130_fd_sc_hd__dfrtp_1 _1131_ (.CLK(clknet_4_0_0_clk),
    .D(_0269_),
    .RESET_B(_0077_),
    .Q(\srfp.register_file[3][13] ));
 sky130_fd_sc_hd__dfrtp_1 _1132_ (.CLK(clknet_4_4_0_clk),
    .D(_0270_),
    .RESET_B(_0078_),
    .Q(\srfp.register_file[3][14] ));
 sky130_fd_sc_hd__dfrtp_2 _1133_ (.CLK(clknet_4_14_0_clk),
    .D(_0271_),
    .RESET_B(_0079_),
    .Q(\srfp.register_file[3][15] ));
 sky130_fd_sc_hd__dfrtp_2 _1134_ (.CLK(clknet_4_9_0_clk),
    .D(_0272_),
    .RESET_B(_0080_),
    .Q(\srfp.register_file[3][16] ));
 sky130_fd_sc_hd__dfrtp_1 _1135_ (.CLK(clknet_4_13_0_clk),
    .D(_0273_),
    .RESET_B(_0081_),
    .Q(\srfp.register_file[3][17] ));
 sky130_fd_sc_hd__dfrtp_1 _1136_ (.CLK(clknet_4_14_0_clk),
    .D(_0274_),
    .RESET_B(_0082_),
    .Q(\srfp.register_file[3][18] ));
 sky130_fd_sc_hd__dfrtp_2 _1137_ (.CLK(clknet_4_10_0_clk),
    .D(_0275_),
    .RESET_B(_0083_),
    .Q(\srfp.register_file[3][19] ));
 sky130_fd_sc_hd__dfrtp_1 _1138_ (.CLK(clknet_4_8_0_clk),
    .D(_0276_),
    .RESET_B(_0084_),
    .Q(\srfp.register_file[3][20] ));
 sky130_fd_sc_hd__dfrtp_1 _1139_ (.CLK(clknet_4_14_0_clk),
    .D(_0277_),
    .RESET_B(_0085_),
    .Q(\srfp.register_file[3][21] ));
 sky130_fd_sc_hd__dfrtp_4 _1140_ (.CLK(clknet_4_9_0_clk),
    .D(_0278_),
    .RESET_B(_0086_),
    .Q(\srfp.register_file[3][22] ));
 sky130_fd_sc_hd__dfrtp_1 _1141_ (.CLK(clknet_4_14_0_clk),
    .D(_0279_),
    .RESET_B(_0087_),
    .Q(\srfp.register_file[3][23] ));
 sky130_fd_sc_hd__dfrtp_4 _1142_ (.CLK(clknet_4_9_0_clk),
    .D(_0280_),
    .RESET_B(_0088_),
    .Q(\srfp.register_file[3][24] ));
 sky130_fd_sc_hd__dfrtp_4 _1143_ (.CLK(clknet_4_9_0_clk),
    .D(_0281_),
    .RESET_B(_0089_),
    .Q(\srfp.register_file[3][25] ));
 sky130_fd_sc_hd__dfrtp_1 _1144_ (.CLK(clknet_4_11_0_clk),
    .D(_0282_),
    .RESET_B(_0090_),
    .Q(\srfp.register_file[3][26] ));
 sky130_fd_sc_hd__dfrtp_1 _1145_ (.CLK(clknet_4_3_0_clk),
    .D(_0283_),
    .RESET_B(_0091_),
    .Q(\srfp.register_file[3][27] ));
 sky130_fd_sc_hd__dfrtp_1 _1146_ (.CLK(clknet_4_11_0_clk),
    .D(_0284_),
    .RESET_B(_0092_),
    .Q(\srfp.register_file[3][28] ));
 sky130_fd_sc_hd__dfrtp_1 _1147_ (.CLK(clknet_4_6_0_clk),
    .D(_0285_),
    .RESET_B(_0093_),
    .Q(\srfp.register_file[3][29] ));
 sky130_fd_sc_hd__dfrtp_1 _1148_ (.CLK(clknet_4_13_0_clk),
    .D(_0286_),
    .RESET_B(_0094_),
    .Q(\srfp.register_file[3][30] ));
 sky130_fd_sc_hd__dfrtp_1 _1149_ (.CLK(clknet_4_4_0_clk),
    .D(_0287_),
    .RESET_B(_0095_),
    .Q(\srfp.register_file[3][31] ));
 sky130_fd_sc_hd__dfrtp_1 _1150_ (.CLK(clknet_4_1_0_clk),
    .D(_0288_),
    .RESET_B(_0096_),
    .Q(\srfp.register_file[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1151_ (.CLK(clknet_4_11_0_clk),
    .D(_0289_),
    .RESET_B(_0097_),
    .Q(\srfp.register_file[2][1] ));
 sky130_fd_sc_hd__dfrtp_2 _1152_ (.CLK(clknet_4_11_0_clk),
    .D(_0290_),
    .RESET_B(_0098_),
    .Q(\srfp.register_file[2][2] ));
 sky130_fd_sc_hd__dfrtp_2 _1153_ (.CLK(clknet_4_3_0_clk),
    .D(_0291_),
    .RESET_B(_0099_),
    .Q(\srfp.register_file[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1154_ (.CLK(clknet_4_8_0_clk),
    .D(_0292_),
    .RESET_B(_0100_),
    .Q(\srfp.register_file[2][4] ));
 sky130_fd_sc_hd__dfrtp_4 _1155_ (.CLK(clknet_4_6_0_clk),
    .D(_0293_),
    .RESET_B(_0101_),
    .Q(\srfp.register_file[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1156_ (.CLK(clknet_4_6_0_clk),
    .D(_0294_),
    .RESET_B(_0102_),
    .Q(\srfp.register_file[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1157_ (.CLK(clknet_4_10_0_clk),
    .D(_0295_),
    .RESET_B(_0103_),
    .Q(\srfp.register_file[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1158_ (.CLK(clknet_4_3_0_clk),
    .D(_0296_),
    .RESET_B(_0104_),
    .Q(\srfp.register_file[2][8] ));
 sky130_fd_sc_hd__dfrtp_1 _1159_ (.CLK(clknet_4_12_0_clk),
    .D(_0297_),
    .RESET_B(_0105_),
    .Q(\srfp.register_file[2][9] ));
 sky130_fd_sc_hd__dfrtp_2 _1160_ (.CLK(clknet_4_8_0_clk),
    .D(_0298_),
    .RESET_B(_0106_),
    .Q(\srfp.register_file[2][10] ));
 sky130_fd_sc_hd__dfrtp_4 _1161_ (.CLK(clknet_4_3_0_clk),
    .D(_0299_),
    .RESET_B(_0107_),
    .Q(\srfp.register_file[2][11] ));
 sky130_fd_sc_hd__dfrtp_1 _1162_ (.CLK(clknet_4_7_0_clk),
    .D(_0300_),
    .RESET_B(_0108_),
    .Q(\srfp.register_file[2][12] ));
 sky130_fd_sc_hd__dfrtp_1 _1163_ (.CLK(clknet_4_0_0_clk),
    .D(_0301_),
    .RESET_B(_0109_),
    .Q(\srfp.register_file[2][13] ));
 sky130_fd_sc_hd__dfrtp_1 _1164_ (.CLK(clknet_4_1_0_clk),
    .D(_0302_),
    .RESET_B(_0110_),
    .Q(\srfp.register_file[2][14] ));
 sky130_fd_sc_hd__dfrtp_2 _1165_ (.CLK(clknet_4_11_0_clk),
    .D(_0303_),
    .RESET_B(_0111_),
    .Q(\srfp.register_file[2][15] ));
 sky130_fd_sc_hd__dfrtp_4 _1166_ (.CLK(clknet_4_15_0_clk),
    .D(_0304_),
    .RESET_B(_0112_),
    .Q(\srfp.register_file[2][16] ));
 sky130_fd_sc_hd__dfrtp_1 _1167_ (.CLK(clknet_4_10_0_clk),
    .D(_0305_),
    .RESET_B(_0113_),
    .Q(\srfp.register_file[2][17] ));
 sky130_fd_sc_hd__dfrtp_1 _1168_ (.CLK(clknet_4_12_0_clk),
    .D(_0306_),
    .RESET_B(_0114_),
    .Q(\srfp.register_file[2][18] ));
 sky130_fd_sc_hd__dfrtp_4 _1169_ (.CLK(clknet_4_12_0_clk),
    .D(_0307_),
    .RESET_B(_0115_),
    .Q(\srfp.register_file[2][19] ));
 sky130_fd_sc_hd__dfrtp_4 _1170_ (.CLK(clknet_4_12_0_clk),
    .D(_0308_),
    .RESET_B(_0116_),
    .Q(\srfp.register_file[2][20] ));
 sky130_fd_sc_hd__dfrtp_1 _1171_ (.CLK(clknet_4_12_0_clk),
    .D(_0309_),
    .RESET_B(_0117_),
    .Q(\srfp.register_file[2][21] ));
 sky130_fd_sc_hd__dfrtp_1 _1172_ (.CLK(clknet_4_6_0_clk),
    .D(_0310_),
    .RESET_B(_0118_),
    .Q(\srfp.register_file[2][22] ));
 sky130_fd_sc_hd__dfrtp_2 _1173_ (.CLK(clknet_4_8_0_clk),
    .D(_0311_),
    .RESET_B(_0119_),
    .Q(\srfp.register_file[2][23] ));
 sky130_fd_sc_hd__dfrtp_4 _1174_ (.CLK(clknet_4_1_0_clk),
    .D(_0312_),
    .RESET_B(_0120_),
    .Q(\srfp.register_file[2][24] ));
 sky130_fd_sc_hd__dfrtp_2 _1175_ (.CLK(clknet_4_2_0_clk),
    .D(_0313_),
    .RESET_B(_0121_),
    .Q(\srfp.register_file[2][25] ));
 sky130_fd_sc_hd__dfrtp_1 _1176_ (.CLK(clknet_4_13_0_clk),
    .D(_0314_),
    .RESET_B(_0122_),
    .Q(\srfp.register_file[2][26] ));
 sky130_fd_sc_hd__dfrtp_1 _1177_ (.CLK(clknet_4_8_0_clk),
    .D(_0315_),
    .RESET_B(_0123_),
    .Q(\srfp.register_file[2][27] ));
 sky130_fd_sc_hd__dfrtp_1 _1178_ (.CLK(clknet_4_10_0_clk),
    .D(_0316_),
    .RESET_B(_0124_),
    .Q(\srfp.register_file[2][28] ));
 sky130_fd_sc_hd__dfrtp_2 _1179_ (.CLK(clknet_4_15_0_clk),
    .D(_0317_),
    .RESET_B(_0125_),
    .Q(\srfp.register_file[2][29] ));
 sky130_fd_sc_hd__dfrtp_1 _1180_ (.CLK(clknet_4_13_0_clk),
    .D(_0318_),
    .RESET_B(_0126_),
    .Q(\srfp.register_file[2][30] ));
 sky130_fd_sc_hd__dfrtp_1 _1181_ (.CLK(clknet_4_0_0_clk),
    .D(_0319_),
    .RESET_B(_0127_),
    .Q(\srfp.register_file[2][31] ));
 sky130_fd_sc_hd__dfrtp_1 _1182_ (.CLK(clknet_4_1_0_clk),
    .D(_0320_),
    .RESET_B(_0128_),
    .Q(\srfp.register_file[1][0] ));
 sky130_fd_sc_hd__dfrtp_2 _1183_ (.CLK(clknet_4_13_0_clk),
    .D(_0321_),
    .RESET_B(_0129_),
    .Q(\srfp.register_file[1][1] ));
 sky130_fd_sc_hd__dfrtp_2 _1184_ (.CLK(clknet_4_14_0_clk),
    .D(_0322_),
    .RESET_B(_0130_),
    .Q(\srfp.register_file[1][2] ));
 sky130_fd_sc_hd__dfrtp_2 _1185_ (.CLK(clknet_4_10_0_clk),
    .D(_0323_),
    .RESET_B(_0131_),
    .Q(\srfp.register_file[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1186_ (.CLK(clknet_4_8_0_clk),
    .D(_0324_),
    .RESET_B(_0132_),
    .Q(\srfp.register_file[1][4] ));
 sky130_fd_sc_hd__dfrtp_2 _1187_ (.CLK(clknet_4_4_0_clk),
    .D(_0325_),
    .RESET_B(_0133_),
    .Q(\srfp.register_file[1][5] ));
 sky130_fd_sc_hd__dfrtp_4 _1188_ (.CLK(clknet_4_6_0_clk),
    .D(_0326_),
    .RESET_B(_0134_),
    .Q(\srfp.register_file[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1189_ (.CLK(clknet_4_2_0_clk),
    .D(_0327_),
    .RESET_B(_0135_),
    .Q(\srfp.register_file[1][7] ));
 sky130_fd_sc_hd__dfrtp_2 _1190_ (.CLK(clknet_4_11_0_clk),
    .D(_0328_),
    .RESET_B(_0136_),
    .Q(\srfp.register_file[1][8] ));
 sky130_fd_sc_hd__dfrtp_1 _1191_ (.CLK(clknet_4_15_0_clk),
    .D(_0329_),
    .RESET_B(_0137_),
    .Q(\srfp.register_file[1][9] ));
 sky130_fd_sc_hd__dfrtp_4 _1192_ (.CLK(clknet_4_0_0_clk),
    .D(_0330_),
    .RESET_B(_0138_),
    .Q(\srfp.register_file[1][10] ));
 sky130_fd_sc_hd__dfrtp_4 _1193_ (.CLK(clknet_4_3_0_clk),
    .D(_0331_),
    .RESET_B(_0139_),
    .Q(\srfp.register_file[1][11] ));
 sky130_fd_sc_hd__dfrtp_4 _1194_ (.CLK(clknet_4_7_0_clk),
    .D(_0332_),
    .RESET_B(_0140_),
    .Q(\srfp.register_file[1][12] ));
 sky130_fd_sc_hd__dfrtp_4 _1195_ (.CLK(clknet_4_3_0_clk),
    .D(_0333_),
    .RESET_B(_0141_),
    .Q(\srfp.register_file[1][13] ));
 sky130_fd_sc_hd__dfrtp_1 _1196_ (.CLK(clknet_4_2_0_clk),
    .D(_0334_),
    .RESET_B(_0142_),
    .Q(\srfp.register_file[1][14] ));
 sky130_fd_sc_hd__dfrtp_1 _1197_ (.CLK(clknet_4_9_0_clk),
    .D(_0335_),
    .RESET_B(_0143_),
    .Q(\srfp.register_file[1][15] ));
 sky130_fd_sc_hd__dfrtp_1 _1198_ (.CLK(clknet_4_5_0_clk),
    .D(_0336_),
    .RESET_B(_0144_),
    .Q(\srfp.register_file[1][16] ));
 sky130_fd_sc_hd__dfrtp_2 _1199_ (.CLK(clknet_4_14_0_clk),
    .D(_0337_),
    .RESET_B(_0145_),
    .Q(\srfp.register_file[1][17] ));
 sky130_fd_sc_hd__dfrtp_1 _1200_ (.CLK(clknet_4_8_0_clk),
    .D(_0338_),
    .RESET_B(_0146_),
    .Q(\srfp.register_file[1][18] ));
 sky130_fd_sc_hd__dfrtp_4 _1201_ (.CLK(clknet_4_0_0_clk),
    .D(_0339_),
    .RESET_B(_0147_),
    .Q(\srfp.register_file[1][19] ));
 sky130_fd_sc_hd__dfrtp_1 _1202_ (.CLK(clknet_4_3_0_clk),
    .D(_0340_),
    .RESET_B(_0148_),
    .Q(\srfp.register_file[1][20] ));
 sky130_fd_sc_hd__dfrtp_1 _1203_ (.CLK(clknet_4_14_0_clk),
    .D(_0341_),
    .RESET_B(_0149_),
    .Q(\srfp.register_file[1][21] ));
 sky130_fd_sc_hd__dfrtp_4 _1204_ (.CLK(clknet_4_1_0_clk),
    .D(_0342_),
    .RESET_B(_0150_),
    .Q(\srfp.register_file[1][22] ));
 sky130_fd_sc_hd__dfrtp_2 _1205_ (.CLK(clknet_4_11_0_clk),
    .D(_0343_),
    .RESET_B(_0151_),
    .Q(\srfp.register_file[1][23] ));
 sky130_fd_sc_hd__dfrtp_1 _1206_ (.CLK(clknet_4_5_0_clk),
    .D(_0344_),
    .RESET_B(_0152_),
    .Q(\srfp.register_file[1][24] ));
 sky130_fd_sc_hd__dfrtp_1 _1207_ (.CLK(clknet_4_11_0_clk),
    .D(_0345_),
    .RESET_B(_0153_),
    .Q(\srfp.register_file[1][25] ));
 sky130_fd_sc_hd__dfrtp_4 _1208_ (.CLK(clknet_4_3_0_clk),
    .D(_0346_),
    .RESET_B(_0154_),
    .Q(\srfp.register_file[1][26] ));
 sky130_fd_sc_hd__dfrtp_1 _1209_ (.CLK(clknet_4_3_0_clk),
    .D(_0347_),
    .RESET_B(_0155_),
    .Q(\srfp.register_file[1][27] ));
 sky130_fd_sc_hd__dfrtp_1 _1210_ (.CLK(clknet_4_11_0_clk),
    .D(_0348_),
    .RESET_B(_0156_),
    .Q(\srfp.register_file[1][28] ));
 sky130_fd_sc_hd__dfrtp_1 _1211_ (.CLK(clknet_4_0_0_clk),
    .D(_0349_),
    .RESET_B(_0157_),
    .Q(\srfp.register_file[1][29] ));
 sky130_fd_sc_hd__dfrtp_1 _1212_ (.CLK(clknet_4_12_0_clk),
    .D(_0350_),
    .RESET_B(_0158_),
    .Q(\srfp.register_file[1][30] ));
 sky130_fd_sc_hd__dfrtp_2 _1213_ (.CLK(clknet_4_10_0_clk),
    .D(_0351_),
    .RESET_B(_0159_),
    .Q(\srfp.register_file[1][31] ));
 sky130_fd_sc_hd__dfrtp_1 _1214_ (.CLK(clknet_4_1_0_clk),
    .D(_0352_),
    .RESET_B(_0160_),
    .Q(\srfp.register_file[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1215_ (.CLK(clknet_4_11_0_clk),
    .D(_0353_),
    .RESET_B(_0161_),
    .Q(\srfp.register_file[0][1] ));
 sky130_fd_sc_hd__dfrtp_4 _1216_ (.CLK(clknet_4_4_0_clk),
    .D(_0354_),
    .RESET_B(_0162_),
    .Q(\srfp.register_file[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1217_ (.CLK(clknet_4_13_0_clk),
    .D(_0355_),
    .RESET_B(_0163_),
    .Q(\srfp.register_file[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1218_ (.CLK(clknet_4_10_0_clk),
    .D(_0356_),
    .RESET_B(_0164_),
    .Q(\srfp.register_file[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1219_ (.CLK(clknet_4_11_0_clk),
    .D(_0357_),
    .RESET_B(_0165_),
    .Q(\srfp.register_file[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1220_ (.CLK(clknet_4_6_0_clk),
    .D(_0358_),
    .RESET_B(_0166_),
    .Q(\srfp.register_file[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1221_ (.CLK(clknet_4_9_0_clk),
    .D(_0359_),
    .RESET_B(_0167_),
    .Q(\srfp.register_file[0][7] ));
 sky130_fd_sc_hd__dfrtp_4 _1222_ (.CLK(clknet_4_3_0_clk),
    .D(_0360_),
    .RESET_B(_0168_),
    .Q(\srfp.register_file[0][8] ));
 sky130_fd_sc_hd__dfrtp_1 _1223_ (.CLK(clknet_4_8_0_clk),
    .D(_0361_),
    .RESET_B(_0169_),
    .Q(\srfp.register_file[0][9] ));
 sky130_fd_sc_hd__dfrtp_1 _1224_ (.CLK(clknet_4_2_0_clk),
    .D(_0362_),
    .RESET_B(_0170_),
    .Q(\srfp.register_file[0][10] ));
 sky130_fd_sc_hd__dfrtp_4 _1225_ (.CLK(clknet_4_15_0_clk),
    .D(_0363_),
    .RESET_B(_0171_),
    .Q(\srfp.register_file[0][11] ));
 sky130_fd_sc_hd__dfrtp_1 _1226_ (.CLK(clknet_4_7_0_clk),
    .D(_0364_),
    .RESET_B(_0172_),
    .Q(\srfp.register_file[0][12] ));
 sky130_fd_sc_hd__dfrtp_4 _1227_ (.CLK(clknet_4_9_0_clk),
    .D(_0365_),
    .RESET_B(_0173_),
    .Q(\srfp.register_file[0][13] ));
 sky130_fd_sc_hd__dfrtp_1 _1228_ (.CLK(clknet_4_0_0_clk),
    .D(_0366_),
    .RESET_B(_0174_),
    .Q(\srfp.register_file[0][14] ));
 sky130_fd_sc_hd__dfrtp_1 _1229_ (.CLK(clknet_4_9_0_clk),
    .D(_0367_),
    .RESET_B(_0175_),
    .Q(\srfp.register_file[0][15] ));
 sky130_fd_sc_hd__dfrtp_1 _1230_ (.CLK(clknet_4_5_0_clk),
    .D(_0368_),
    .RESET_B(_0176_),
    .Q(\srfp.register_file[0][16] ));
 sky130_fd_sc_hd__dfrtp_1 _1231_ (.CLK(clknet_4_14_0_clk),
    .D(_0369_),
    .RESET_B(_0177_),
    .Q(\srfp.register_file[0][17] ));
 sky130_fd_sc_hd__dfrtp_4 _1232_ (.CLK(clknet_4_12_0_clk),
    .D(_0370_),
    .RESET_B(_0178_),
    .Q(\srfp.register_file[0][18] ));
 sky130_fd_sc_hd__dfrtp_1 _1233_ (.CLK(clknet_4_4_0_clk),
    .D(_0371_),
    .RESET_B(_0179_),
    .Q(\srfp.register_file[0][19] ));
 sky130_fd_sc_hd__dfrtp_1 _1234_ (.CLK(clknet_4_5_0_clk),
    .D(_0372_),
    .RESET_B(_0180_),
    .Q(\srfp.register_file[0][20] ));
 sky130_fd_sc_hd__dfrtp_1 _1235_ (.CLK(clknet_4_11_0_clk),
    .D(_0373_),
    .RESET_B(_0181_),
    .Q(\srfp.register_file[0][21] ));
 sky130_fd_sc_hd__dfrtp_1 _1236_ (.CLK(clknet_4_5_0_clk),
    .D(_0374_),
    .RESET_B(_0182_),
    .Q(\srfp.register_file[0][22] ));
 sky130_fd_sc_hd__dfrtp_1 _1237_ (.CLK(clknet_4_15_0_clk),
    .D(_0375_),
    .RESET_B(_0183_),
    .Q(\srfp.register_file[0][23] ));
 sky130_fd_sc_hd__dfrtp_4 _1238_ (.CLK(clknet_4_4_0_clk),
    .D(_0376_),
    .RESET_B(_0184_),
    .Q(\srfp.register_file[0][24] ));
 sky130_fd_sc_hd__dfrtp_1 _1239_ (.CLK(clknet_4_12_0_clk),
    .D(_0377_),
    .RESET_B(_0185_),
    .Q(\srfp.register_file[0][25] ));
 sky130_fd_sc_hd__dfrtp_1 _1240_ (.CLK(clknet_4_13_0_clk),
    .D(_0378_),
    .RESET_B(_0186_),
    .Q(\srfp.register_file[0][26] ));
 sky130_fd_sc_hd__dfrtp_1 _1241_ (.CLK(clknet_4_10_0_clk),
    .D(_0379_),
    .RESET_B(_0187_),
    .Q(\srfp.register_file[0][27] ));
 sky130_fd_sc_hd__dfrtp_1 _1242_ (.CLK(clknet_4_2_0_clk),
    .D(_0380_),
    .RESET_B(_0188_),
    .Q(\srfp.register_file[0][28] ));
 sky130_fd_sc_hd__dfrtp_1 _1243_ (.CLK(clknet_4_4_0_clk),
    .D(_0381_),
    .RESET_B(_0189_),
    .Q(\srfp.register_file[0][29] ));
 sky130_fd_sc_hd__dfrtp_1 _1244_ (.CLK(clknet_4_14_0_clk),
    .D(_0382_),
    .RESET_B(_0190_),
    .Q(\srfp.register_file[0][30] ));
 sky130_fd_sc_hd__dfrtp_1 _1245_ (.CLK(clknet_4_1_0_clk),
    .D(_0383_),
    .RESET_B(_0191_),
    .Q(\srfp.register_file[0][31] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_8 fanout100 (.A(_0389_),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 fanout101 (.A(_0389_),
    .X(net101));
 sky130_fd_sc_hd__buf_6 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_6 fanout103 (.A(_0389_),
    .X(net103));
 sky130_fd_sc_hd__buf_6 fanout104 (.A(net107),
    .X(net104));
 sky130_fd_sc_hd__buf_6 fanout105 (.A(net107),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_8 fanout107 (.A(_0388_),
    .X(net107));
 sky130_fd_sc_hd__buf_6 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_4 fanout109 (.A(_0387_),
    .X(net109));
 sky130_fd_sc_hd__buf_6 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__buf_6 fanout111 (.A(_0387_),
    .X(net111));
 sky130_fd_sc_hd__buf_6 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(_0386_),
    .X(net113));
 sky130_fd_sc_hd__buf_6 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_6 fanout115 (.A(_0386_),
    .X(net115));
 sky130_fd_sc_hd__buf_6 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_8 fanout117 (.A(net119),
    .X(net117));
 sky130_fd_sc_hd__buf_6 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_8 fanout119 (.A(_0385_),
    .X(net119));
 sky130_fd_sc_hd__buf_6 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__buf_6 fanout121 (.A(net123),
    .X(net121));
 sky130_fd_sc_hd__buf_6 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__buf_6 fanout123 (.A(_0384_),
    .X(net123));
 sky130_fd_sc_hd__buf_6 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_8 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_8 fanout126 (.A(net130),
    .X(net126));
 sky130_fd_sc_hd__buf_6 fanout127 (.A(net129),
    .X(net127));
 sky130_fd_sc_hd__buf_6 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_8 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_6 fanout130 (.A(net135),
    .X(net130));
 sky130_fd_sc_hd__buf_6 fanout131 (.A(net135),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net135),
    .X(net132));
 sky130_fd_sc_hd__buf_8 fanout133 (.A(net135),
    .X(net133));
 sky130_fd_sc_hd__buf_6 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_6 fanout135 (.A(net4),
    .X(net135));
 sky130_fd_sc_hd__buf_6 fanout136 (.A(net145),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(net145),
    .X(net137));
 sky130_fd_sc_hd__buf_6 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net145),
    .X(net139));
 sky130_fd_sc_hd__buf_6 fanout140 (.A(net145),
    .X(net140));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net145),
    .X(net141));
 sky130_fd_sc_hd__buf_6 fanout142 (.A(net144),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_4 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net4),
    .X(net145));
 sky130_fd_sc_hd__buf_8 fanout146 (.A(net149),
    .X(net146));
 sky130_fd_sc_hd__buf_8 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_8 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_8 fanout149 (.A(net4),
    .X(net149));
 sky130_fd_sc_hd__buf_8 fanout150 (.A(net3),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 fanout151 (.A(net3),
    .X(net151));
 sky130_fd_sc_hd__buf_6 fanout152 (.A(net2),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(net2),
    .X(net153));
 sky130_fd_sc_hd__buf_6 fanout154 (.A(net1),
    .X(net154));
 sky130_fd_sc_hd__buf_4 fanout73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(_0398_),
    .X(net74));
 sky130_fd_sc_hd__buf_4 fanout75 (.A(_0398_),
    .X(net75));
 sky130_fd_sc_hd__buf_2 fanout76 (.A(_0398_),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(_0397_),
    .X(net78));
 sky130_fd_sc_hd__buf_4 fanout79 (.A(_0397_),
    .X(net79));
 sky130_fd_sc_hd__buf_2 fanout80 (.A(_0397_),
    .X(net80));
 sky130_fd_sc_hd__buf_6 fanout81 (.A(net83),
    .X(net81));
 sky130_fd_sc_hd__buf_6 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_4 fanout83 (.A(_0396_),
    .X(net83));
 sky130_fd_sc_hd__buf_6 fanout84 (.A(_0394_),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(_0394_),
    .X(net85));
 sky130_fd_sc_hd__buf_6 fanout86 (.A(_0394_),
    .X(net86));
 sky130_fd_sc_hd__buf_4 fanout87 (.A(_0394_),
    .X(net87));
 sky130_fd_sc_hd__buf_4 fanout88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 fanout89 (.A(_0393_),
    .X(net89));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(_0393_),
    .X(net90));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(_0393_),
    .X(net91));
 sky130_fd_sc_hd__buf_4 fanout92 (.A(_0392_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 fanout93 (.A(_0392_),
    .X(net93));
 sky130_fd_sc_hd__buf_6 fanout94 (.A(_0392_),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(_0392_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_8 fanout96 (.A(_0390_),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 fanout97 (.A(_0390_),
    .X(net97));
 sky130_fd_sc_hd__buf_4 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(_0390_),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(read_address[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(write_data[11]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(write_data[12]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(write_data[13]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(write_data[14]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(write_data[15]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(write_data[16]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(write_data[17]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(write_data[18]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(write_data[19]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(write_data[1]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(read_address[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input20 (.A(write_data[20]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(write_data[21]),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input22 (.A(write_data[22]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(write_data[23]),
    .X(net23));
 sky130_fd_sc_hd__buf_6 input24 (.A(write_data[24]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(write_data[25]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(write_data[26]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(write_data[27]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(write_data[28]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(write_data[29]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(read_address[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(write_data[2]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(write_data[30]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(write_data[31]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(write_data[3]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(write_data[4]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(write_data[5]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(write_data[6]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(write_data[7]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(write_data[8]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(write_data[9]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input4 (.A(reset),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input40 (.A(write_enable),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(write_address[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(write_address[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(write_address[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(write_data[0]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(write_data[10]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 output41 (.A(net41),
    .X(read_data[0]));
 sky130_fd_sc_hd__clkbuf_2 output42 (.A(net42),
    .X(read_data[10]));
 sky130_fd_sc_hd__clkbuf_2 output43 (.A(net43),
    .X(read_data[11]));
 sky130_fd_sc_hd__clkbuf_2 output44 (.A(net44),
    .X(read_data[12]));
 sky130_fd_sc_hd__clkbuf_2 output45 (.A(net45),
    .X(read_data[13]));
 sky130_fd_sc_hd__clkbuf_2 output46 (.A(net46),
    .X(read_data[14]));
 sky130_fd_sc_hd__clkbuf_2 output47 (.A(net47),
    .X(read_data[15]));
 sky130_fd_sc_hd__clkbuf_2 output48 (.A(net48),
    .X(read_data[16]));
 sky130_fd_sc_hd__clkbuf_2 output49 (.A(net49),
    .X(read_data[17]));
 sky130_fd_sc_hd__clkbuf_2 output50 (.A(net50),
    .X(read_data[18]));
 sky130_fd_sc_hd__clkbuf_2 output51 (.A(net51),
    .X(read_data[19]));
 sky130_fd_sc_hd__clkbuf_2 output52 (.A(net52),
    .X(read_data[1]));
 sky130_fd_sc_hd__clkbuf_2 output53 (.A(net53),
    .X(read_data[20]));
 sky130_fd_sc_hd__clkbuf_2 output54 (.A(net54),
    .X(read_data[21]));
 sky130_fd_sc_hd__clkbuf_2 output55 (.A(net55),
    .X(read_data[22]));
 sky130_fd_sc_hd__clkbuf_2 output56 (.A(net56),
    .X(read_data[23]));
 sky130_fd_sc_hd__clkbuf_2 output57 (.A(net57),
    .X(read_data[24]));
 sky130_fd_sc_hd__clkbuf_2 output58 (.A(net58),
    .X(read_data[25]));
 sky130_fd_sc_hd__clkbuf_2 output59 (.A(net59),
    .X(read_data[26]));
 sky130_fd_sc_hd__clkbuf_2 output60 (.A(net60),
    .X(read_data[27]));
 sky130_fd_sc_hd__clkbuf_2 output61 (.A(net61),
    .X(read_data[28]));
 sky130_fd_sc_hd__clkbuf_2 output62 (.A(net62),
    .X(read_data[29]));
 sky130_fd_sc_hd__clkbuf_2 output63 (.A(net63),
    .X(read_data[2]));
 sky130_fd_sc_hd__clkbuf_2 output64 (.A(net64),
    .X(read_data[30]));
 sky130_fd_sc_hd__clkbuf_2 output65 (.A(net65),
    .X(read_data[31]));
 sky130_fd_sc_hd__clkbuf_2 output66 (.A(net66),
    .X(read_data[3]));
 sky130_fd_sc_hd__clkbuf_2 output67 (.A(net67),
    .X(read_data[4]));
 sky130_fd_sc_hd__clkbuf_2 output68 (.A(net68),
    .X(read_data[5]));
 sky130_fd_sc_hd__clkbuf_2 output69 (.A(net69),
    .X(read_data[6]));
 sky130_fd_sc_hd__clkbuf_2 output70 (.A(net70),
    .X(read_data[7]));
 sky130_fd_sc_hd__clkbuf_2 output71 (.A(net71),
    .X(read_data[8]));
 sky130_fd_sc_hd__clkbuf_2 output72 (.A(net72),
    .X(read_data[9]));
endmodule

