//Filepaths added by humans
`include "../../Dpath/sim/queue.v"
`include "../../Dpath/sim/Counter.v"
`include "../../Dpath/sim/Decoder.v"
`include "../../RegisterFiles/sim/VectorRegFile.v"
`include "../../Dpath/sim/ALU.v"
`include "../../RegisterFiles/sim/Scalar_Register_File.v"
`include "../../RegisterFiles/sim/Predicate_Register_File.v"
module TopModule (
    input logic clk,
    input logic reset,

    // Receive interface for load_queue
    input logic [63:0] load_recv_msg,
    input logic load_recv_val,
    output logic load_recv_rdy,

    // Receive interface for instruction_queue
    input logic [31:0] instruction_recv_msg,
    input logic instruction_recv_val,
    output logic instruction_recv_rdy,

    // Send interface for store_queue
    output logic [31:0] store_send_msg,
    output logic store_send_val,
    input logic store_send_rdy
);

    // Internal signals for send interface of load_queue and instruction_queue
    logic [63:0] load_send_msg;
    logic load_send_val;
    logic load_send_rdy;

    logic [31:0] instruction_send_msg;
    logic instruction_send_val;
    logic instruction_send_rdy;

    // Internal signals for receive interface of store_queue
    logic [31:0] store_recv_msg;
    logic store_recv_val;
    logic store_recv_rdy;

    // Internal signals for Decoder
    logic clock_enable;
    logic clock_bypass;
    logic [4:0] vector_reg_write_select;
    logic [4:0] reg_file_addr1;
    logic [4:0] reg_file_addr2;
    logic mux_bit;
    logic vector_reg_write_bit;
    logic predicate_reg_write_bit;
    logic scalar_reg_write_bit;
    logic vector_reg_load_mux_bit;
    logic scalar_reg_load_mux_bit;
    logic [2:0] functional_unit_mux_bit;
    logic add_subtract_bit;
    logic load_store_bit;
    logic [1:0] bitwise_op_select;
    logic [3:0] predicate_op_select;

    // Internal signals for VectorRegFile
    logic [31:0] wb_addr;
    logic [31:0] wb_data;
    logic [31:0] rData1;
    logic [31:0] rData2;

    // New wire for functional_unit_output_mux
    logic [31:0] functional_unit_output_mux;

    // Mux output for VectorRegFile wData
    logic [31:0] wData_mux_out;

    // Mux outputs for VectorRegFile wAddr1 and wAddr2
    logic [4:0] wAddr1_mux_out;
    logic [4:0] wAddr2_mux_out;

    // 2-input muxes for VectorRegFile rAddr1_1 and rAddr2_1
    logic [4:0] rAddr1_1_mux_out;
    logic [4:0] rAddr2_1_mux_out;

    // Internal signals for Scalar_Register_File
    logic [4:0] scalar_read_address;
    logic [4:0] scalar_write_address;
    logic [31:0] scalar_write_data;
    logic scalar_write_enable;
    logic [31:0] scalar_read_data;

    // New signal declaration for vector_write_enable
    logic vector_write_enable;

    // Assign the expression to the new signal
    assign vector_write_enable = (vector_reg_write_bit & !load_store_bit & pred_data_out) | (vector_reg_write_bit & load_store_bit & (wb_addr <= addr_cutoff));

    // New signal declaration for addr_cutoff
    logic [31:0] addr_cutoff;
    assign addr_cutoff = 32'h000003FF;  // Updated to 32'h00000400

    // Modified assignment for scalar_write_address
    assign scalar_write_address = wb_addr[4:0] - addr_cutoff[4:0] - 1;  // Removed -1

    // Modified assignment for scalar_read_address
    assign scalar_read_address = load_store_bit ? scalar_write_address : reg_file_addr2;

    // Conditional assignment for store_recv_msg
    assign store_recv_msg = (wb_addr > addr_cutoff) ? scalar_read_data : rData1;

    // Corrected line
    assign store_recv_val = load_store_bit & !vector_reg_write_bit;

    // Corrected line
    assign load_send_rdy = load_store_bit;

    // Instantiate load_queue
    queue #(.WIDTH(64), .DEPTH(16)) load_queue (
        .clk(clk),
        .reset(reset),
        .recv_msg(load_recv_msg),
        .recv_val(load_recv_val),
        .recv_rdy(load_recv_rdy),
        .send_msg(load_send_msg),
        .send_val(load_send_val),
        .send_rdy(load_send_rdy)
    );

    // Instantiate instruction_queue
    queue #(.WIDTH(32), .DEPTH(16)) instruction_queue (
        .clk(clk),
        .reset(reset),
        .recv_msg(instruction_recv_msg),
        .recv_val(instruction_recv_val),
        .recv_rdy(instruction_recv_rdy),
        .send_msg(instruction_send_msg),
        .send_val(instruction_send_val),
        .send_rdy(instruction_send_rdy)
    );

    // Instantiate store_queue
    queue #(.WIDTH(32), .DEPTH(16)) store_queue (
        .clk(clk),
        .reset(reset),
        .recv_msg(store_recv_msg),
        .recv_val(store_recv_val),
        .recv_rdy(store_recv_rdy),
        .send_msg(store_send_msg),
        .send_val(store_send_val),
        .send_rdy(store_send_rdy)
    );

    // Instantiate Decoder
    Decoder decoder (
        .instruction(instruction_send_msg),
        .instruction_valid(instruction_send_val),
        .reg_file_addr1(reg_file_addr1),
        .reg_file_addr2(reg_file_addr2),
        .mux_bit(mux_bit),
        .vector_reg_write_bit(vector_reg_write_bit),
        .predicate_reg_write_bit(predicate_reg_write_bit),
        .scalar_reg_write_bit(scalar_reg_write_bit),
        .vector_reg_load_mux_bit(vector_reg_load_mux_bit),
        .scalar_reg_load_mux_bit(scalar_reg_load_mux_bit),
        .functional_unit_mux_bit(functional_unit_mux_bit),
        .add_subtract_bit(add_subtract_bit),
        .load_store_bit(load_store_bit),
        .clock_enable(clock_enable),
        .clock_bypass(clock_bypass),
        .bitwise_op_select(bitwise_op_select),
        .predicate_op_select(predicate_op_select),
        .vector_reg_write_select(vector_reg_write_select)
    );

    // Internal signal for Counter
    logic [4:0] counter;
    logic done;

    // Instantiate Counter
    Counter #(.WIDTH(5), .COUNTER_MAX(2**5-1)) counter_module (
        .clk(clk),
        .enable(clock_enable),
        .reset(reset),
        .counter(counter),
        .done(done)
    );

    // OR the done output with clock_bypass and connect this result to instruction_send_rdy
    assign instruction_send_rdy = done | clock_bypass;  // Updated to done | clock_bypass

    // Create new wires for wb_addr and wb_data
    assign wb_addr = load_send_msg[63:32];
    assign wb_data = load_send_msg[31:0];

    // 2-input mux for VectorRegFile wData
    assign wData_mux_out = load_store_bit ? wb_data : functional_unit_output_mux;

    // 2-input muxes for VectorRegFile wAddr1 and wAddr2
    assign wAddr1_mux_out = load_store_bit ? wb_addr[9:5] : vector_reg_write_select;
    assign wAddr2_mux_out = load_store_bit ? wb_addr[4:0] : counter;

    // 2-input muxes for VectorRegFile rAddr1_1 and rAddr2_1
    assign rAddr1_1_mux_out = load_store_bit ? wb_addr[9:5] : reg_file_addr1;
    assign rAddr2_1_mux_out = load_store_bit ? wb_addr[4:0] : counter;

    // Instantiate VectorRegFile
    VectorRegFile #(.ADDR_WIDTH(5), .DATA_WIDTH(32), .NUM_REG(32), .NUM_ELE(32)) reg_file (
        .clk(clk),
        .reset(reset),
        .rAddr1_1(rAddr1_1_mux_out),
        .rAddr2_1(rAddr2_1_mux_out),
        .rData1(rData1),
        .rAddr1_2(reg_file_addr2),
        .rAddr2_2(counter),
        .rData2(rData2),
        .wAddr1(wAddr1_mux_out),
        .wAddr2(wAddr2_mux_out),
        .wData(wData_mux_out),
        .wEnable(vector_write_enable)  // Updated to use the new signal
    );

    // Instantiate ALU
    ALU #(32) alu (
        .A(rData1),
        .B(rData2),  // Updated input
        .C(scalar_read_data),  // Updated input
        .AddSub(add_subtract_bit),
        .muxControl(mux_bit),
        .outputControl(functional_unit_mux_bit),
        .bitwiseControl(bitwise_op_select),
        .compControl(predicate_op_select),
        .finalResult(functional_unit_output_mux),
        .predicate(pred_data_in) // Updated input
    );

    // Assignments for Scalar_Register_File
    assign scalar_write_data = wb_data;
    assign scalar_write_enable = load_store_bit & vector_reg_write_bit & (wb_addr > addr_cutoff);

    // Instantiate Scalar_Register_File
    Scalar_Register_File #(
        .REG_DEPTH(32),
        .REG_WIDTH(32),
        .ADDR_WIDTH(5)
    ) scalar_reg_file (
        .clk(clk),
        .reset(reset),  // Added reset connection
        .read_address(scalar_read_address),
        .write_address(scalar_write_address),
        .write_data(scalar_write_data),
        .write_enable(scalar_write_enable),
        .read_data(scalar_read_data)
    );

    // Internal signals for Predicate_Register_File
    logic [4:0] pred_read_addr1, pred_read_addr2;
    logic [4:0] pred_write_addr1, pred_write_addr2;
    logic pred_write_enable;
    logic pred_data_out;
    logic pred_data_in;

    // Assignments for Predicate_Register_File
    assign pred_read_addr1 = vector_reg_write_select; // Updated line
    assign pred_read_addr2 = counter;
    assign pred_write_addr1 = vector_reg_write_select;
    assign pred_write_addr2 = counter;
    assign pred_write_enable = predicate_reg_write_bit;

    // Instantiate Predicate_Register_File
    Predicate_Register_File #(
        .ADDR_WIDTH(5),
        .DATA_WIDTH(1),
        .NUM_REGISTERS(32)
    ) predicate_reg_file (
        .clk(clk),
        .reset(reset),
        .read_addr1(pred_read_addr1),
        .read_addr2(pred_read_addr2),
        .write_addr1(pred_write_addr1),
        .write_addr2(pred_write_addr2),
        .write_enable(pred_write_enable),
        .data_out(pred_data_out),
        .data_in(pred_data_in)
    );

endmodule
