magic
tech sky130A
magscale 1 2
timestamp 1692313518
<< viali >>
rect 3157 26537 3191 26571
rect 8033 26537 8067 26571
rect 27353 26537 27387 26571
rect 29929 26537 29963 26571
rect 32505 26537 32539 26571
rect 35081 26537 35115 26571
rect 37657 26537 37691 26571
rect 6929 26469 6963 26503
rect 20361 26469 20395 26503
rect 38485 26469 38519 26503
rect 2329 26401 2363 26435
rect 4261 26401 4295 26435
rect 13277 26401 13311 26435
rect 18337 26401 18371 26435
rect 25605 26401 25639 26435
rect 29193 26401 29227 26435
rect 36553 26401 36587 26435
rect 2053 26333 2087 26367
rect 3985 26333 4019 26367
rect 6653 26333 6687 26367
rect 9137 26333 9171 26367
rect 11713 26333 11747 26367
rect 13001 26333 13035 26367
rect 14933 26333 14967 26367
rect 17141 26333 17175 26367
rect 18153 26333 18187 26367
rect 20177 26333 20211 26367
rect 22017 26333 22051 26367
rect 23305 26333 23339 26367
rect 25329 26333 25363 26367
rect 27261 26333 27295 26367
rect 28457 26333 28491 26367
rect 28595 26333 28629 26367
rect 28733 26333 28767 26367
rect 29837 26333 29871 26367
rect 30757 26333 30791 26367
rect 34989 26333 35023 26367
rect 36277 26333 36311 26367
rect 38301 26333 38335 26367
rect 3065 26265 3099 26299
rect 7941 26265 7975 26299
rect 9413 26265 9447 26299
rect 15209 26265 15243 26299
rect 16957 26265 16991 26299
rect 23581 26265 23615 26299
rect 31125 26265 31159 26299
rect 32413 26265 32447 26299
rect 37565 26265 37599 26299
rect 38025 26265 38059 26299
rect 11897 26197 11931 26231
rect 22201 26197 22235 26231
rect 1777 25993 1811 26027
rect 18061 25993 18095 26027
rect 38301 25925 38335 25959
rect 1685 25857 1719 25891
rect 13185 25857 13219 25891
rect 16129 25857 16163 25891
rect 16865 25857 16899 25891
rect 17969 25857 18003 25891
rect 29377 25857 29411 25891
rect 37565 25857 37599 25891
rect 18245 25789 18279 25823
rect 13277 25653 13311 25687
rect 16221 25653 16255 25687
rect 17049 25653 17083 25687
rect 17601 25653 17635 25687
rect 29377 25653 29411 25687
rect 37657 25653 37691 25687
rect 38393 25653 38427 25687
rect 1777 25449 1811 25483
rect 36645 25449 36679 25483
rect 29837 25381 29871 25415
rect 38669 25381 38703 25415
rect 7481 25313 7515 25347
rect 15669 25313 15703 25347
rect 18245 25313 18279 25347
rect 27169 25313 27203 25347
rect 30389 25313 30423 25347
rect 1685 25245 1719 25279
rect 15393 25245 15427 25279
rect 18061 25245 18095 25279
rect 26893 25245 26927 25279
rect 32689 25245 32723 25279
rect 36185 25245 36219 25279
rect 36553 25245 36587 25279
rect 36737 25245 36771 25279
rect 38485 25245 38519 25279
rect 13093 25177 13127 25211
rect 30205 25177 30239 25211
rect 33057 25177 33091 25211
rect 6837 25109 6871 25143
rect 7205 25109 7239 25143
rect 7297 25109 7331 25143
rect 13369 25109 13403 25143
rect 17141 25109 17175 25143
rect 28641 25109 28675 25143
rect 30297 25109 30331 25143
rect 36369 25109 36403 25143
rect 13001 24837 13035 24871
rect 17601 24837 17635 24871
rect 23581 24837 23615 24871
rect 32597 24837 32631 24871
rect 34805 24837 34839 24871
rect 36185 24837 36219 24871
rect 36737 24837 36771 24871
rect 14013 24769 14047 24803
rect 14841 24769 14875 24803
rect 18153 24769 18187 24803
rect 25145 24769 25179 24803
rect 30297 24769 30331 24803
rect 35173 24769 35207 24803
rect 35265 24769 35299 24803
rect 35357 24769 35391 24803
rect 36553 24769 36587 24803
rect 36645 24769 36679 24803
rect 38025 24769 38059 24803
rect 13093 24701 13127 24735
rect 13277 24701 13311 24735
rect 15025 24701 15059 24735
rect 18061 24701 18095 24735
rect 23673 24701 23707 24735
rect 23857 24701 23891 24735
rect 32321 24701 32355 24735
rect 34713 24701 34747 24735
rect 36093 24701 36127 24735
rect 38301 24701 38335 24735
rect 17601 24633 17635 24667
rect 24961 24633 24995 24667
rect 12633 24565 12667 24599
rect 14105 24565 14139 24599
rect 18337 24565 18371 24599
rect 23213 24565 23247 24599
rect 30113 24565 30147 24599
rect 34069 24565 34103 24599
rect 8309 24361 8343 24395
rect 15853 24361 15887 24395
rect 16221 24361 16255 24395
rect 17877 24361 17911 24395
rect 28181 24361 28215 24395
rect 35449 24361 35483 24395
rect 36829 24361 36863 24395
rect 12633 24293 12667 24327
rect 6193 24225 6227 24259
rect 13185 24225 13219 24259
rect 14841 24225 14875 24259
rect 18337 24225 18371 24259
rect 18521 24225 18555 24259
rect 26801 24225 26835 24259
rect 34989 24225 35023 24259
rect 35541 24225 35575 24259
rect 1685 24157 1719 24191
rect 5917 24157 5951 24191
rect 8217 24157 8251 24191
rect 15853 24157 15887 24191
rect 16037 24157 16071 24191
rect 26893 24157 26927 24191
rect 27077 24157 27111 24191
rect 28089 24157 28123 24191
rect 31861 24157 31895 24191
rect 32597 24157 32631 24191
rect 35081 24157 35115 24191
rect 36461 24157 36495 24191
rect 36553 24157 36587 24191
rect 36921 24157 36955 24191
rect 2237 24089 2271 24123
rect 9321 24089 9355 24123
rect 18245 24089 18279 24123
rect 27537 24089 27571 24123
rect 32965 24089 32999 24123
rect 7665 24021 7699 24055
rect 9413 24021 9447 24055
rect 13001 24021 13035 24055
rect 13093 24021 13127 24055
rect 14289 24021 14323 24055
rect 14657 24021 14691 24055
rect 14749 24021 14783 24055
rect 31953 24021 31987 24055
rect 35817 24021 35851 24055
rect 37105 24021 37139 24055
rect 5089 23817 5123 23851
rect 8217 23817 8251 23851
rect 13645 23817 13679 23851
rect 14105 23817 14139 23851
rect 4997 23681 5031 23715
rect 6929 23681 6963 23715
rect 7021 23681 7055 23715
rect 9137 23681 9171 23715
rect 13001 23681 13035 23715
rect 14013 23681 14047 23715
rect 14841 23681 14875 23715
rect 16957 23681 16991 23715
rect 17417 23681 17451 23715
rect 17693 23681 17727 23715
rect 24869 23681 24903 23715
rect 32689 23681 32723 23715
rect 32781 23681 32815 23715
rect 34897 23681 34931 23715
rect 34989 23681 35023 23715
rect 35357 23681 35391 23715
rect 7205 23613 7239 23647
rect 8309 23613 8343 23647
rect 8401 23613 8435 23647
rect 9413 23613 9447 23647
rect 14197 23613 14231 23647
rect 15025 23613 15059 23647
rect 25145 23613 25179 23647
rect 32873 23613 32907 23647
rect 6561 23477 6595 23511
rect 7849 23477 7883 23511
rect 13093 23477 13127 23511
rect 18245 23477 18279 23511
rect 26617 23477 26651 23511
rect 32321 23477 32355 23511
rect 35357 23477 35391 23511
rect 35541 23477 35575 23511
rect 9321 23273 9355 23307
rect 9505 23273 9539 23307
rect 25605 23273 25639 23307
rect 31861 23273 31895 23307
rect 6837 23137 6871 23171
rect 7021 23137 7055 23171
rect 13553 23137 13587 23171
rect 23949 23137 23983 23171
rect 2237 23069 2271 23103
rect 2881 23069 2915 23103
rect 10701 23069 10735 23103
rect 14289 23069 14323 23103
rect 23673 23069 23707 23103
rect 25513 23069 25547 23103
rect 2329 23001 2363 23035
rect 9137 23001 9171 23035
rect 11253 23001 11287 23035
rect 31677 23001 31711 23035
rect 2973 22933 3007 22967
rect 6377 22933 6411 22967
rect 6745 22933 6779 22967
rect 9337 22933 9371 22967
rect 13001 22933 13035 22967
rect 13369 22933 13403 22967
rect 13461 22933 13495 22967
rect 14381 22933 14415 22967
rect 23305 22933 23339 22967
rect 23765 22933 23799 22967
rect 31877 22933 31911 22967
rect 32045 22933 32079 22967
rect 2237 22729 2271 22763
rect 4747 22729 4781 22763
rect 21281 22729 21315 22763
rect 31769 22729 31803 22763
rect 1685 22661 1719 22695
rect 4537 22661 4571 22695
rect 10425 22661 10459 22695
rect 14197 22661 14231 22695
rect 32321 22661 32355 22695
rect 3617 22593 3651 22627
rect 5733 22593 5767 22627
rect 5825 22593 5859 22627
rect 10241 22593 10275 22627
rect 10701 22593 10735 22627
rect 12909 22593 12943 22627
rect 13921 22593 13955 22627
rect 18429 22593 18463 22627
rect 24317 22593 24351 22627
rect 24409 22593 24443 22627
rect 31401 22593 31435 22627
rect 31585 22593 31619 22627
rect 13093 22525 13127 22559
rect 15945 22525 15979 22559
rect 18705 22525 18739 22559
rect 19533 22525 19567 22559
rect 19809 22525 19843 22559
rect 24593 22525 24627 22559
rect 33057 22525 33091 22559
rect 23949 22457 23983 22491
rect 1777 22389 1811 22423
rect 3709 22389 3743 22423
rect 4721 22389 4755 22423
rect 4905 22389 4939 22423
rect 6009 22389 6043 22423
rect 31585 22389 31619 22423
rect 3341 22049 3375 22083
rect 4629 22049 4663 22083
rect 10701 22049 10735 22083
rect 13553 22049 13587 22083
rect 14933 22049 14967 22083
rect 16589 22049 16623 22083
rect 31585 22049 31619 22083
rect 32965 22049 32999 22083
rect 14841 21981 14875 22015
rect 15853 21981 15887 22015
rect 16497 21981 16531 22015
rect 18613 21981 18647 22015
rect 28549 21981 28583 22015
rect 30205 21981 30239 22015
rect 31309 21981 31343 22015
rect 10977 21913 11011 21947
rect 13277 21913 13311 21947
rect 15945 21913 15979 21947
rect 2697 21845 2731 21879
rect 3065 21845 3099 21879
rect 3157 21845 3191 21879
rect 3985 21845 4019 21879
rect 4353 21845 4387 21879
rect 4445 21845 4479 21879
rect 12449 21845 12483 21879
rect 12909 21845 12943 21879
rect 13369 21845 13403 21879
rect 18705 21845 18739 21879
rect 28641 21845 28675 21879
rect 30297 21845 30331 21879
rect 32413 21845 32447 21879
rect 32781 21845 32815 21879
rect 32873 21845 32907 21879
rect 4077 21641 4111 21675
rect 13185 21641 13219 21675
rect 26525 21641 26559 21675
rect 12909 21573 12943 21607
rect 17233 21573 17267 21607
rect 31217 21573 31251 21607
rect 3985 21505 4019 21539
rect 12633 21505 12667 21539
rect 12817 21505 12851 21539
rect 13025 21505 13059 21539
rect 24777 21505 24811 21539
rect 28273 21505 28307 21539
rect 35725 21505 35759 21539
rect 16957 21437 16991 21471
rect 25053 21437 25087 21471
rect 28549 21437 28583 21471
rect 31309 21437 31343 21471
rect 31493 21437 31527 21471
rect 35817 21369 35851 21403
rect 18705 21301 18739 21335
rect 30021 21301 30055 21335
rect 30849 21301 30883 21335
rect 27813 21097 27847 21131
rect 29929 21097 29963 21131
rect 11161 20961 11195 20995
rect 25145 20961 25179 20995
rect 25421 20961 25455 20995
rect 28365 20961 28399 20995
rect 36921 20961 36955 20995
rect 1593 20893 1627 20927
rect 3985 20893 4019 20927
rect 12449 20893 12483 20927
rect 13277 20893 13311 20927
rect 13737 20893 13771 20927
rect 31033 20893 31067 20927
rect 34897 20893 34931 20927
rect 1869 20825 1903 20859
rect 11069 20825 11103 20859
rect 12909 20825 12943 20859
rect 29745 20825 29779 20859
rect 35173 20825 35207 20859
rect 38485 20825 38519 20859
rect 38669 20825 38703 20859
rect 4077 20757 4111 20791
rect 10609 20757 10643 20791
rect 10977 20757 11011 20791
rect 26893 20757 26927 20791
rect 28181 20757 28215 20791
rect 28273 20757 28307 20791
rect 29945 20757 29979 20791
rect 30113 20757 30147 20791
rect 31125 20757 31159 20791
rect 27537 20553 27571 20587
rect 28733 20553 28767 20587
rect 33149 20553 33183 20587
rect 36185 20553 36219 20587
rect 4629 20485 4663 20519
rect 12127 20485 12161 20519
rect 29193 20485 29227 20519
rect 33609 20485 33643 20519
rect 4537 20417 4571 20451
rect 11713 20417 11747 20451
rect 21189 20417 21223 20451
rect 22017 20417 22051 20451
rect 22753 20417 22787 20451
rect 23673 20417 23707 20451
rect 29101 20417 29135 20451
rect 33517 20417 33551 20451
rect 36093 20417 36127 20451
rect 2237 20349 2271 20383
rect 2513 20349 2547 20383
rect 27629 20349 27663 20383
rect 27721 20349 27755 20383
rect 29377 20349 29411 20383
rect 33793 20349 33827 20383
rect 12265 20281 12299 20315
rect 22201 20281 22235 20315
rect 3985 20213 4019 20247
rect 12081 20213 12115 20247
rect 21373 20213 21407 20247
rect 22845 20213 22879 20247
rect 23765 20213 23799 20247
rect 27169 20213 27203 20247
rect 6009 20009 6043 20043
rect 14473 20009 14507 20043
rect 33057 20009 33091 20043
rect 22845 19941 22879 19975
rect 5825 19873 5859 19907
rect 13737 19873 13771 19907
rect 18521 19873 18555 19907
rect 21005 19873 21039 19907
rect 21097 19873 21131 19907
rect 2697 19805 2731 19839
rect 6009 19805 6043 19839
rect 12449 19805 12483 19839
rect 12817 19805 12851 19839
rect 13185 19805 13219 19839
rect 18705 19805 18739 19839
rect 19451 19805 19485 19839
rect 19717 19805 19751 19839
rect 20637 19805 20671 19839
rect 21649 19805 21683 19839
rect 21833 19805 21867 19839
rect 22017 19805 22051 19839
rect 22661 19805 22695 19839
rect 31309 19805 31343 19839
rect 5457 19737 5491 19771
rect 5733 19737 5767 19771
rect 14381 19737 14415 19771
rect 20545 19737 20579 19771
rect 21925 19737 21959 19771
rect 31585 19737 31619 19771
rect 2789 19669 2823 19703
rect 6193 19669 6227 19703
rect 18889 19669 18923 19703
rect 22201 19669 22235 19703
rect 15301 19465 15335 19499
rect 20111 19465 20145 19499
rect 26341 19465 26375 19499
rect 31309 19465 31343 19499
rect 36093 19465 36127 19499
rect 36461 19465 36495 19499
rect 4445 19397 4479 19431
rect 5641 19397 5675 19431
rect 14933 19397 14967 19431
rect 15025 19397 15059 19431
rect 19901 19397 19935 19431
rect 31033 19397 31067 19431
rect 35449 19397 35483 19431
rect 35541 19397 35575 19431
rect 4353 19329 4387 19363
rect 5457 19329 5491 19363
rect 5733 19329 5767 19363
rect 5825 19329 5859 19363
rect 11897 19329 11931 19363
rect 12449 19329 12483 19363
rect 14749 19329 14783 19363
rect 15117 19329 15151 19363
rect 17509 19329 17543 19363
rect 17601 19329 17635 19363
rect 20821 19329 20855 19363
rect 22385 19329 22419 19363
rect 24593 19329 24627 19363
rect 30757 19329 30791 19363
rect 30941 19329 30975 19363
rect 31125 19329 31159 19363
rect 35265 19329 35299 19363
rect 36553 19329 36587 19363
rect 12725 19261 12759 19295
rect 21373 19261 21407 19295
rect 22661 19261 22695 19295
rect 24869 19261 24903 19295
rect 36645 19261 36679 19295
rect 6009 19193 6043 19227
rect 14197 19193 14231 19227
rect 11897 19125 11931 19159
rect 20085 19125 20119 19159
rect 20269 19125 20303 19159
rect 24133 19125 24167 19159
rect 34989 19125 35023 19159
rect 28273 18921 28307 18955
rect 27077 18853 27111 18887
rect 30665 18853 30699 18887
rect 20821 18785 20855 18819
rect 23673 18785 23707 18819
rect 26249 18785 26283 18819
rect 26341 18785 26375 18819
rect 26433 18785 26467 18819
rect 27537 18785 27571 18819
rect 32321 18785 32355 18819
rect 32597 18785 32631 18819
rect 34345 18785 34379 18819
rect 37473 18785 37507 18819
rect 1685 18717 1719 18751
rect 5641 18717 5675 18751
rect 6285 18717 6319 18751
rect 12081 18717 12115 18751
rect 19901 18717 19935 18751
rect 23489 18717 23523 18751
rect 24961 18717 24995 18751
rect 28181 18717 28215 18751
rect 35725 18717 35759 18751
rect 37197 18717 37231 18751
rect 6377 18649 6411 18683
rect 17785 18649 17819 18683
rect 18521 18649 18555 18683
rect 20177 18649 20211 18683
rect 21097 18649 21131 18683
rect 25421 18649 25455 18683
rect 27629 18649 27663 18683
rect 30941 18649 30975 18683
rect 31217 18649 31251 18683
rect 36461 18649 36495 18683
rect 1777 18581 1811 18615
rect 5733 18581 5767 18615
rect 12173 18581 12207 18615
rect 22569 18581 22603 18615
rect 23029 18581 23063 18615
rect 23397 18581 23431 18615
rect 26065 18581 26099 18615
rect 27537 18581 27571 18615
rect 31125 18581 31159 18615
rect 20637 18377 20671 18411
rect 21281 18377 21315 18411
rect 24041 18377 24075 18411
rect 24593 18377 24627 18411
rect 25053 18377 25087 18411
rect 26525 18377 26559 18411
rect 31309 18377 31343 18411
rect 37565 18377 37599 18411
rect 2973 18309 3007 18343
rect 17509 18309 17543 18343
rect 19809 18309 19843 18343
rect 19901 18309 19935 18343
rect 31217 18309 31251 18343
rect 13185 18241 13219 18275
rect 17325 18241 17359 18275
rect 17601 18241 17635 18275
rect 17693 18241 17727 18275
rect 19625 18241 19659 18275
rect 19993 18241 20027 18275
rect 20913 18241 20947 18275
rect 21373 18241 21407 18275
rect 22569 18241 22603 18275
rect 23949 18241 23983 18275
rect 24961 18241 24995 18275
rect 25881 18241 25915 18275
rect 26617 18241 26651 18275
rect 27169 18241 27203 18275
rect 35633 18241 35667 18275
rect 37473 18241 37507 18275
rect 2697 18173 2731 18207
rect 4445 18173 4479 18207
rect 13461 18173 13495 18207
rect 23305 18173 23339 18207
rect 25145 18173 25179 18207
rect 26341 18173 26375 18207
rect 27353 18173 27387 18207
rect 31401 18173 31435 18207
rect 36461 18173 36495 18207
rect 20177 18105 20211 18139
rect 21097 18105 21131 18139
rect 14933 18037 14967 18071
rect 17877 18037 17911 18071
rect 21005 18037 21039 18071
rect 26157 18037 26191 18071
rect 26249 18037 26283 18071
rect 30849 18037 30883 18071
rect 25973 17833 26007 17867
rect 26157 17833 26191 17867
rect 21097 17765 21131 17799
rect 24593 17765 24627 17799
rect 26709 17765 26743 17799
rect 15945 17697 15979 17731
rect 21741 17697 21775 17731
rect 22293 17697 22327 17731
rect 22569 17697 22603 17731
rect 25237 17697 25271 17731
rect 31033 17697 31067 17731
rect 31309 17697 31343 17731
rect 33057 17697 33091 17731
rect 2053 17629 2087 17663
rect 2697 17629 2731 17663
rect 15669 17629 15703 17663
rect 20269 17629 20303 17663
rect 24961 17629 24995 17663
rect 27169 17629 27203 17663
rect 29745 17629 29779 17663
rect 33793 17629 33827 17663
rect 21557 17561 21591 17595
rect 25053 17561 25087 17595
rect 25789 17561 25823 17595
rect 25989 17561 26023 17595
rect 26709 17561 26743 17595
rect 2145 17493 2179 17527
rect 2789 17493 2823 17527
rect 17417 17493 17451 17527
rect 20361 17493 20395 17527
rect 21465 17493 21499 17527
rect 24041 17493 24075 17527
rect 27261 17493 27295 17527
rect 27445 17493 27479 17527
rect 29837 17493 29871 17527
rect 33885 17493 33919 17527
rect 7665 17289 7699 17323
rect 23949 17289 23983 17323
rect 26433 17289 26467 17323
rect 30113 17289 30147 17323
rect 32965 17289 32999 17323
rect 5273 17221 5307 17255
rect 14381 17221 14415 17255
rect 17141 17221 17175 17255
rect 23213 17221 23247 17255
rect 25237 17221 25271 17255
rect 27261 17221 27295 17255
rect 31585 17221 31619 17255
rect 32597 17221 32631 17255
rect 32689 17221 32723 17255
rect 34253 17221 34287 17255
rect 35449 17221 35483 17255
rect 1593 17153 1627 17187
rect 5181 17153 5215 17187
rect 8033 17153 8067 17187
rect 14105 17153 14139 17187
rect 16865 17153 16899 17187
rect 22569 17153 22603 17187
rect 23857 17153 23891 17187
rect 24501 17153 24535 17187
rect 25881 17153 25915 17187
rect 26065 17153 26099 17187
rect 26157 17153 26191 17187
rect 26249 17153 26283 17187
rect 30021 17153 30055 17187
rect 30849 17153 30883 17187
rect 32321 17153 32355 17187
rect 32414 17153 32448 17187
rect 32827 17153 32861 17187
rect 34161 17153 34195 17187
rect 35081 17153 35115 17187
rect 38485 17153 38519 17187
rect 2605 17085 2639 17119
rect 2881 17085 2915 17119
rect 5365 17085 5399 17119
rect 8125 17085 8159 17119
rect 8217 17085 8251 17119
rect 16129 17085 16163 17119
rect 18889 17085 18923 17119
rect 19349 17085 19383 17119
rect 19625 17085 19659 17119
rect 30297 17085 30331 17119
rect 34345 17085 34379 17119
rect 33793 17017 33827 17051
rect 38669 17017 38703 17051
rect 1685 16949 1719 16983
rect 4353 16949 4387 16983
rect 4813 16949 4847 16983
rect 21097 16949 21131 16983
rect 27353 16949 27387 16983
rect 29653 16949 29687 16983
rect 1961 16745 1995 16779
rect 12817 16745 12851 16779
rect 26617 16745 26651 16779
rect 13001 16677 13035 16711
rect 33057 16677 33091 16711
rect 33149 16677 33183 16711
rect 35449 16677 35483 16711
rect 4813 16609 4847 16643
rect 4905 16609 4939 16643
rect 21005 16609 21039 16643
rect 21281 16609 21315 16643
rect 23673 16609 23707 16643
rect 23765 16609 23799 16643
rect 25329 16609 25363 16643
rect 30665 16609 30699 16643
rect 30757 16609 30791 16643
rect 32781 16609 32815 16643
rect 2605 16541 2639 16575
rect 3249 16541 3283 16575
rect 5549 16541 5583 16575
rect 6193 16541 6227 16575
rect 13553 16541 13587 16575
rect 13645 16541 13679 16575
rect 14657 16541 14691 16575
rect 14933 16541 14967 16575
rect 15025 16541 15059 16575
rect 15761 16541 15795 16575
rect 17233 16541 17267 16575
rect 17325 16541 17359 16575
rect 17877 16541 17911 16575
rect 26617 16541 26651 16575
rect 27353 16541 27387 16575
rect 31401 16541 31435 16575
rect 33241 16541 33275 16575
rect 33517 16541 33551 16575
rect 34161 16541 34195 16575
rect 34897 16541 34931 16575
rect 35265 16541 35299 16575
rect 35909 16541 35943 16575
rect 36553 16541 36587 16575
rect 12863 16507 12897 16541
rect 1685 16473 1719 16507
rect 12633 16473 12667 16507
rect 14841 16473 14875 16507
rect 16313 16473 16347 16507
rect 24593 16473 24627 16507
rect 27629 16473 27663 16507
rect 32229 16473 32263 16507
rect 34253 16473 34287 16507
rect 35081 16473 35115 16507
rect 35173 16473 35207 16507
rect 2697 16405 2731 16439
rect 3341 16405 3375 16439
rect 4353 16405 4387 16439
rect 4721 16405 4755 16439
rect 5641 16405 5675 16439
rect 6285 16405 6319 16439
rect 15209 16405 15243 16439
rect 17969 16405 18003 16439
rect 22753 16405 22787 16439
rect 23213 16405 23247 16439
rect 23581 16405 23615 16439
rect 29101 16405 29135 16439
rect 30205 16405 30239 16439
rect 30573 16405 30607 16439
rect 33425 16405 33459 16439
rect 36001 16405 36035 16439
rect 36645 16405 36679 16439
rect 11805 16201 11839 16235
rect 23765 16201 23799 16235
rect 29193 16201 29227 16235
rect 5641 16133 5675 16167
rect 8953 16133 8987 16167
rect 9137 16133 9171 16167
rect 12449 16133 12483 16167
rect 13553 16133 13587 16167
rect 17141 16133 17175 16167
rect 22293 16133 22327 16167
rect 29929 16133 29963 16167
rect 33425 16133 33459 16167
rect 1593 16065 1627 16099
rect 5089 16065 5123 16099
rect 10977 16065 11011 16099
rect 11713 16065 11747 16099
rect 13277 16065 13311 16099
rect 15853 16065 15887 16099
rect 16037 16065 16071 16099
rect 16129 16065 16163 16099
rect 16865 16065 16899 16099
rect 27445 16065 27479 16099
rect 32505 16065 32539 16099
rect 33149 16065 33183 16099
rect 35817 16065 35851 16099
rect 36645 16065 36679 16099
rect 37473 16065 37507 16099
rect 2237 15997 2271 16031
rect 2513 15997 2547 16031
rect 9229 15997 9263 16031
rect 15025 15997 15059 16031
rect 16313 15997 16347 16031
rect 22017 15997 22051 16031
rect 27721 15997 27755 16031
rect 29653 15997 29687 16031
rect 35909 15997 35943 16031
rect 36001 15997 36035 16031
rect 8677 15929 8711 15963
rect 11069 15929 11103 15963
rect 12725 15929 12759 15963
rect 15577 15929 15611 15963
rect 15945 15929 15979 15963
rect 1685 15861 1719 15895
rect 3985 15861 4019 15895
rect 31401 15861 31435 15895
rect 32597 15861 32631 15895
rect 34897 15861 34931 15895
rect 35449 15861 35483 15895
rect 36737 15861 36771 15895
rect 37565 15861 37599 15895
rect 2697 15657 2731 15691
rect 5733 15657 5767 15691
rect 8217 15657 8251 15691
rect 10044 15657 10078 15691
rect 13737 15657 13771 15691
rect 26433 15657 26467 15691
rect 28457 15657 28491 15691
rect 33885 15657 33919 15691
rect 34069 15657 34103 15691
rect 19809 15589 19843 15623
rect 25237 15589 25271 15623
rect 28089 15589 28123 15623
rect 32781 15589 32815 15623
rect 32873 15589 32907 15623
rect 3157 15521 3191 15555
rect 3341 15521 3375 15555
rect 9229 15521 9263 15555
rect 9781 15521 9815 15555
rect 11989 15521 12023 15555
rect 15945 15521 15979 15555
rect 16221 15521 16255 15555
rect 22845 15521 22879 15555
rect 25697 15521 25731 15555
rect 28917 15521 28951 15555
rect 29009 15521 29043 15555
rect 30205 15521 30239 15555
rect 35081 15521 35115 15555
rect 38117 15521 38151 15555
rect 1593 15453 1627 15487
rect 3985 15453 4019 15487
rect 6193 15453 6227 15487
rect 6837 15453 6871 15487
rect 8125 15453 8159 15487
rect 9137 15453 9171 15487
rect 18153 15453 18187 15487
rect 19533 15453 19567 15487
rect 21097 15453 21131 15487
rect 23857 15453 23891 15487
rect 26341 15453 26375 15487
rect 28825 15453 28859 15487
rect 29929 15453 29963 15487
rect 31401 15453 31435 15487
rect 31677 15453 31711 15487
rect 31769 15453 31803 15487
rect 32965 15453 32999 15487
rect 33057 15453 33091 15487
rect 33241 15453 33275 15487
rect 37933 15453 37967 15487
rect 1869 15385 1903 15419
rect 4261 15385 4295 15419
rect 6285 15385 6319 15419
rect 12265 15385 12299 15419
rect 14289 15385 14323 15419
rect 15025 15385 15059 15419
rect 21373 15385 21407 15419
rect 25789 15385 25823 15419
rect 31585 15385 31619 15419
rect 32505 15385 32539 15419
rect 33701 15385 33735 15419
rect 35357 15385 35391 15419
rect 37105 15385 37139 15419
rect 38025 15385 38059 15419
rect 3065 15317 3099 15351
rect 6929 15317 6963 15351
rect 11529 15317 11563 15351
rect 17693 15317 17727 15351
rect 18337 15317 18371 15351
rect 23949 15317 23983 15351
rect 24869 15317 24903 15351
rect 25697 15317 25731 15351
rect 31953 15317 31987 15351
rect 33901 15317 33935 15351
rect 37565 15317 37599 15351
rect 7113 15113 7147 15147
rect 7941 15113 7975 15147
rect 10333 15113 10367 15147
rect 11069 15113 11103 15147
rect 11713 15113 11747 15147
rect 12173 15113 12207 15147
rect 17417 15113 17451 15147
rect 18153 15113 18187 15147
rect 18521 15113 18555 15147
rect 21097 15113 21131 15147
rect 28833 15113 28867 15147
rect 31217 15113 31251 15147
rect 37841 15113 37875 15147
rect 3249 15045 3283 15079
rect 5549 15045 5583 15079
rect 5733 15045 5767 15079
rect 5825 15045 5859 15079
rect 6837 15045 6871 15079
rect 13369 15045 13403 15079
rect 14105 15045 14139 15079
rect 16957 15045 16991 15079
rect 18613 15045 18647 15079
rect 19533 15045 19567 15079
rect 19625 15045 19659 15079
rect 23397 15045 23431 15079
rect 30849 15045 30883 15079
rect 31065 15045 31099 15079
rect 35173 15045 35207 15079
rect 38485 15045 38519 15079
rect 2237 14977 2271 15011
rect 6561 14977 6595 15011
rect 6745 14977 6779 15011
rect 6929 14977 6963 15011
rect 7573 14977 7607 15011
rect 7757 14977 7791 15011
rect 10977 14977 11011 15011
rect 12081 14977 12115 15011
rect 15485 14977 15519 15011
rect 19349 14977 19383 15011
rect 19717 14977 19751 15011
rect 21189 14977 21223 15011
rect 22017 14977 22051 15011
rect 23121 14977 23155 15011
rect 28273 14977 28307 15011
rect 28457 14977 28491 15011
rect 28549 14977 28583 15011
rect 28646 14977 28680 15011
rect 29377 14977 29411 15011
rect 32321 14977 32355 15011
rect 34897 14977 34931 15011
rect 37749 14977 37783 15011
rect 38669 14977 38703 15011
rect 2053 14909 2087 14943
rect 2973 14909 3007 14943
rect 8585 14909 8619 14943
rect 8861 14909 8895 14943
rect 12265 14909 12299 14943
rect 16129 14909 16163 14943
rect 17509 14909 17543 14943
rect 18705 14909 18739 14943
rect 21373 14909 21407 14943
rect 22201 14909 22235 14943
rect 25145 14909 25179 14943
rect 29929 14909 29963 14943
rect 32597 14909 32631 14943
rect 5273 14841 5307 14875
rect 16957 14841 16991 14875
rect 2421 14773 2455 14807
rect 4721 14773 4755 14807
rect 7757 14773 7791 14807
rect 17693 14773 17727 14807
rect 19901 14773 19935 14807
rect 20729 14773 20763 14807
rect 31033 14773 31067 14807
rect 34069 14773 34103 14807
rect 36645 14773 36679 14807
rect 1777 14569 1811 14603
rect 2145 14569 2179 14603
rect 2697 14569 2731 14603
rect 4169 14569 4203 14603
rect 10333 14569 10367 14603
rect 19625 14569 19659 14603
rect 38025 14569 38059 14603
rect 13737 14501 13771 14535
rect 22569 14501 22603 14535
rect 37381 14501 37415 14535
rect 3157 14433 3191 14467
rect 3341 14433 3375 14467
rect 4997 14433 5031 14467
rect 9597 14433 9631 14467
rect 9781 14433 9815 14467
rect 10885 14433 10919 14467
rect 16221 14433 16255 14467
rect 20269 14433 20303 14467
rect 25053 14433 25087 14467
rect 28917 14433 28951 14467
rect 29009 14433 29043 14467
rect 30297 14433 30331 14467
rect 31033 14433 31067 14467
rect 34989 14433 35023 14467
rect 1869 14365 1903 14399
rect 1961 14365 1995 14399
rect 7205 14365 7239 14399
rect 11805 14365 11839 14399
rect 13093 14365 13127 14399
rect 13241 14365 13275 14399
rect 13599 14365 13633 14399
rect 14841 14365 14875 14399
rect 15945 14365 15979 14399
rect 18429 14365 18463 14399
rect 19993 14365 20027 14399
rect 20821 14365 20855 14399
rect 27813 14365 27847 14399
rect 33425 14365 33459 14399
rect 33793 14365 33827 14399
rect 37197 14365 37231 14399
rect 37933 14365 37967 14399
rect 1685 14297 1719 14331
rect 3065 14297 3099 14331
rect 3985 14297 4019 14331
rect 4201 14297 4235 14331
rect 5273 14297 5307 14331
rect 7941 14297 7975 14331
rect 10701 14297 10735 14331
rect 12265 14297 12299 14331
rect 13369 14297 13403 14331
rect 13461 14297 13495 14331
rect 15393 14297 15427 14331
rect 17969 14297 18003 14331
rect 18705 14297 18739 14331
rect 21097 14297 21131 14331
rect 25329 14297 25363 14331
rect 27905 14297 27939 14331
rect 28825 14297 28859 14331
rect 30113 14297 30147 14331
rect 31309 14297 31343 14331
rect 35265 14297 35299 14331
rect 4353 14229 4387 14263
rect 6745 14229 6779 14263
rect 9137 14229 9171 14263
rect 9505 14229 9539 14263
rect 10793 14229 10827 14263
rect 20085 14229 20119 14263
rect 26801 14229 26835 14263
rect 28457 14229 28491 14263
rect 29745 14229 29779 14263
rect 30205 14229 30239 14263
rect 32781 14229 32815 14263
rect 36737 14229 36771 14263
rect 8309 14025 8343 14059
rect 8677 14025 8711 14059
rect 10793 14025 10827 14059
rect 29929 14025 29963 14059
rect 32321 14025 32355 14059
rect 34161 14025 34195 14059
rect 34713 14025 34747 14059
rect 35449 14025 35483 14059
rect 35817 14025 35851 14059
rect 2053 13957 2087 13991
rect 10425 13957 10459 13991
rect 10641 13957 10675 13991
rect 16221 13957 16255 13991
rect 19717 13957 19751 13991
rect 21465 13957 21499 13991
rect 28457 13957 28491 13991
rect 33793 13957 33827 13991
rect 37565 13957 37599 13991
rect 4077 13889 4111 13923
rect 6929 13889 6963 13923
rect 8769 13889 8803 13923
rect 9505 13889 9539 13923
rect 11989 13889 12023 13923
rect 12725 13889 12759 13923
rect 15301 13889 15335 13923
rect 15393 13889 15427 13923
rect 16129 13889 16163 13923
rect 17233 13889 17267 13923
rect 18613 13889 18647 13923
rect 22201 13889 22235 13923
rect 24869 13889 24903 13923
rect 27169 13889 27203 13923
rect 28181 13889 28215 13923
rect 30573 13889 30607 13923
rect 31309 13889 31343 13923
rect 32689 13889 32723 13923
rect 33609 13889 33643 13923
rect 33885 13889 33919 13923
rect 33977 13889 34011 13923
rect 34621 13889 34655 13923
rect 36737 13889 36771 13923
rect 37473 13889 37507 13923
rect 38117 13889 38151 13923
rect 1777 13821 1811 13855
rect 3525 13821 3559 13855
rect 5825 13821 5859 13855
rect 7757 13821 7791 13855
rect 8861 13821 8895 13855
rect 9781 13821 9815 13855
rect 14473 13821 14507 13855
rect 15577 13821 15611 13855
rect 17325 13821 17359 13855
rect 17417 13821 17451 13855
rect 19165 13821 19199 13855
rect 23949 13821 23983 13855
rect 27261 13821 27295 13855
rect 30665 13821 30699 13855
rect 32781 13821 32815 13855
rect 32965 13821 32999 13855
rect 35909 13821 35943 13855
rect 36001 13821 36035 13855
rect 36829 13821 36863 13855
rect 14933 13753 14967 13787
rect 4334 13685 4368 13719
rect 10609 13685 10643 13719
rect 12081 13685 12115 13719
rect 12988 13685 13022 13719
rect 16865 13685 16899 13719
rect 22464 13685 22498 13719
rect 25132 13685 25166 13719
rect 26617 13685 26651 13719
rect 31401 13685 31435 13719
rect 38209 13685 38243 13719
rect 3985 13481 4019 13515
rect 8309 13481 8343 13515
rect 8493 13481 8527 13515
rect 14749 13481 14783 13515
rect 16037 13481 16071 13515
rect 18429 13481 18463 13515
rect 18797 13481 18831 13515
rect 23121 13481 23155 13515
rect 24961 13481 24995 13515
rect 32321 13481 32355 13515
rect 36645 13481 36679 13515
rect 16313 13413 16347 13447
rect 18291 13413 18325 13447
rect 23305 13413 23339 13447
rect 27353 13413 27387 13447
rect 34069 13413 34103 13447
rect 4537 13345 4571 13379
rect 5917 13345 5951 13379
rect 10793 13345 10827 13379
rect 15301 13345 15335 13379
rect 18521 13345 18555 13379
rect 20453 13345 20487 13379
rect 25605 13345 25639 13379
rect 26617 13345 26651 13379
rect 26801 13345 26835 13379
rect 27997 13345 28031 13379
rect 30573 13345 30607 13379
rect 33333 13345 33367 13379
rect 34897 13345 34931 13379
rect 2605 13277 2639 13311
rect 3249 13277 3283 13311
rect 3341 13277 3375 13311
rect 5181 13277 5215 13311
rect 9689 13277 9723 13311
rect 10333 13277 10367 13311
rect 12909 13277 12943 13311
rect 13185 13277 13219 13311
rect 13461 13277 13495 13311
rect 13553 13277 13587 13311
rect 16405 13277 16439 13311
rect 16497 13277 16531 13311
rect 16773 13277 16807 13311
rect 17233 13277 17267 13311
rect 19441 13277 19475 13311
rect 19625 13277 19659 13311
rect 19809 13277 19843 13311
rect 22477 13277 22511 13311
rect 23857 13277 23891 13311
rect 25421 13277 25455 13311
rect 27813 13277 27847 13311
rect 28549 13277 28583 13311
rect 29745 13277 29779 13311
rect 33149 13277 33183 13311
rect 33977 13277 34011 13311
rect 37565 13277 37599 13311
rect 1685 13209 1719 13243
rect 4353 13209 4387 13243
rect 6193 13209 6227 13243
rect 8125 13209 8159 13243
rect 9781 13209 9815 13243
rect 11069 13209 11103 13243
rect 13369 13209 13403 13243
rect 15209 13209 15243 13243
rect 17509 13209 17543 13243
rect 18153 13209 18187 13243
rect 19717 13209 19751 13243
rect 20729 13209 20763 13243
rect 22937 13209 22971 13243
rect 25329 13209 25363 13243
rect 27721 13209 27755 13243
rect 29837 13209 29871 13243
rect 30849 13209 30883 13243
rect 35173 13209 35207 13243
rect 38301 13209 38335 13243
rect 1777 13141 1811 13175
rect 2697 13141 2731 13175
rect 4445 13141 4479 13175
rect 5273 13141 5307 13175
rect 7665 13141 7699 13175
rect 8325 13141 8359 13175
rect 10425 13141 10459 13175
rect 12541 13141 12575 13175
rect 13737 13141 13771 13175
rect 15117 13141 15151 13175
rect 16681 13141 16715 13175
rect 19993 13141 20027 13175
rect 23137 13141 23171 13175
rect 23949 13141 23983 13175
rect 26157 13141 26191 13175
rect 26525 13141 26559 13175
rect 28641 13141 28675 13175
rect 32781 13141 32815 13175
rect 33241 13141 33275 13175
rect 37657 13141 37691 13175
rect 38393 13141 38427 13175
rect 7573 12937 7607 12971
rect 7941 12937 7975 12971
rect 8033 12937 8067 12971
rect 11713 12937 11747 12971
rect 13553 12937 13587 12971
rect 14749 12937 14783 12971
rect 16145 12937 16179 12971
rect 18613 12937 18647 12971
rect 25237 12937 25271 12971
rect 25881 12937 25915 12971
rect 26341 12937 26375 12971
rect 31493 12937 31527 12971
rect 2513 12869 2547 12903
rect 4261 12869 4295 12903
rect 9781 12869 9815 12903
rect 13185 12869 13219 12903
rect 13385 12869 13419 12903
rect 15971 12869 16005 12903
rect 17141 12869 17175 12903
rect 27997 12869 28031 12903
rect 28917 12869 28951 12903
rect 29009 12869 29043 12903
rect 30021 12869 30055 12903
rect 32965 12869 32999 12903
rect 34897 12869 34931 12903
rect 1593 12801 1627 12835
rect 5181 12801 5215 12835
rect 5825 12801 5859 12835
rect 6929 12801 6963 12835
rect 8769 12801 8803 12835
rect 9689 12801 9723 12835
rect 10333 12801 10367 12835
rect 10977 12801 11011 12835
rect 12081 12801 12115 12835
rect 12173 12801 12207 12835
rect 14013 12801 14047 12835
rect 14105 12801 14139 12835
rect 15301 12801 15335 12835
rect 16865 12801 16899 12835
rect 19073 12801 19107 12835
rect 22017 12801 22051 12835
rect 22937 12801 22971 12835
rect 25145 12801 25179 12835
rect 26249 12801 26283 12835
rect 27537 12801 27571 12835
rect 28733 12801 28767 12835
rect 29101 12801 29135 12835
rect 29745 12801 29779 12835
rect 32781 12801 32815 12835
rect 33057 12801 33091 12835
rect 33149 12801 33183 12835
rect 33793 12801 33827 12835
rect 34805 12801 34839 12835
rect 35725 12801 35759 12835
rect 37565 12801 37599 12835
rect 38209 12801 38243 12835
rect 2237 12733 2271 12767
rect 5917 12733 5951 12767
rect 8217 12733 8251 12767
rect 8953 12733 8987 12767
rect 12357 12733 12391 12767
rect 15209 12733 15243 12767
rect 15485 12733 15519 12767
rect 19349 12733 19383 12767
rect 21097 12733 21131 12767
rect 22201 12733 22235 12767
rect 23213 12733 23247 12767
rect 26525 12733 26559 12767
rect 34989 12733 35023 12767
rect 36001 12733 36035 12767
rect 10425 12665 10459 12699
rect 15025 12665 15059 12699
rect 16313 12665 16347 12699
rect 37657 12665 37691 12699
rect 1685 12597 1719 12631
rect 5273 12597 5307 12631
rect 7021 12597 7055 12631
rect 11069 12597 11103 12631
rect 13369 12597 13403 12631
rect 15117 12597 15151 12631
rect 16129 12597 16163 12631
rect 24685 12597 24719 12631
rect 29285 12597 29319 12631
rect 33333 12597 33367 12631
rect 33885 12597 33919 12631
rect 34437 12597 34471 12631
rect 38301 12597 38335 12631
rect 12541 12393 12575 12427
rect 13737 12393 13771 12427
rect 15485 12393 15519 12427
rect 16037 12393 16071 12427
rect 17785 12393 17819 12427
rect 20361 12393 20395 12427
rect 21281 12393 21315 12427
rect 32597 12393 32631 12427
rect 35081 12393 35115 12427
rect 36001 12393 36035 12427
rect 37933 12393 37967 12427
rect 5733 12325 5767 12359
rect 9781 12325 9815 12359
rect 11069 12325 11103 12359
rect 12725 12325 12759 12359
rect 20250 12325 20284 12359
rect 32781 12325 32815 12359
rect 36829 12325 36863 12359
rect 7481 12257 7515 12291
rect 16497 12257 16531 12291
rect 16681 12257 16715 12291
rect 18613 12257 18647 12291
rect 20453 12257 20487 12291
rect 20821 12257 20855 12291
rect 21833 12257 21867 12291
rect 25697 12257 25731 12291
rect 28549 12257 28583 12291
rect 30205 12257 30239 12291
rect 30481 12257 30515 12291
rect 31953 12257 31987 12291
rect 33793 12257 33827 12291
rect 1961 12189 1995 12223
rect 2605 12189 2639 12223
rect 3249 12189 3283 12223
rect 3985 12189 4019 12223
rect 6285 12189 6319 12223
rect 8401 12189 8435 12223
rect 9689 12189 9723 12223
rect 10333 12189 10367 12223
rect 11529 12189 11563 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 13553 12189 13587 12223
rect 14289 12189 14323 12223
rect 14933 12189 14967 12223
rect 15301 12189 15335 12223
rect 17233 12189 17267 12223
rect 17509 12189 17543 12223
rect 17601 12189 17635 12223
rect 18429 12189 18463 12223
rect 19441 12189 19475 12223
rect 20085 12189 20119 12223
rect 22477 12189 22511 12223
rect 23857 12189 23891 12223
rect 24869 12189 24903 12223
rect 28273 12189 28307 12223
rect 35817 12189 35851 12223
rect 35909 12189 35943 12223
rect 36737 12189 36771 12223
rect 37841 12189 37875 12223
rect 38485 12189 38519 12223
rect 2053 12121 2087 12155
rect 4261 12121 4295 12155
rect 7389 12121 7423 12155
rect 11069 12121 11103 12155
rect 12357 12121 12391 12155
rect 12573 12121 12607 12155
rect 13461 12121 13495 12155
rect 15117 12121 15151 12155
rect 15209 12121 15243 12155
rect 17417 12121 17451 12155
rect 19533 12121 19567 12155
rect 21741 12121 21775 12155
rect 22753 12121 22787 12155
rect 25973 12121 26007 12155
rect 32413 12121 32447 12155
rect 33609 12121 33643 12155
rect 33701 12121 33735 12155
rect 34989 12121 35023 12155
rect 38577 12121 38611 12155
rect 2697 12053 2731 12087
rect 3341 12053 3375 12087
rect 6377 12053 6411 12087
rect 6929 12053 6963 12087
rect 7297 12053 7331 12087
rect 8493 12053 8527 12087
rect 10425 12053 10459 12087
rect 11621 12053 11655 12087
rect 11805 12053 11839 12087
rect 14381 12053 14415 12087
rect 16405 12053 16439 12087
rect 21649 12053 21683 12087
rect 23949 12053 23983 12087
rect 24961 12053 24995 12087
rect 27445 12053 27479 12087
rect 27905 12053 27939 12087
rect 28365 12053 28399 12087
rect 32613 12053 32647 12087
rect 33241 12053 33275 12087
rect 36185 12053 36219 12087
rect 6561 11849 6595 11883
rect 7205 11849 7239 11883
rect 16313 11849 16347 11883
rect 19533 11849 19567 11883
rect 20085 11849 20119 11883
rect 20453 11849 20487 11883
rect 20545 11849 20579 11883
rect 25329 11849 25363 11883
rect 28917 11849 28951 11883
rect 31125 11849 31159 11883
rect 32689 11849 32723 11883
rect 33057 11849 33091 11883
rect 36645 11849 36679 11883
rect 13185 11781 13219 11815
rect 17509 11781 17543 11815
rect 22293 11781 22327 11815
rect 25697 11781 25731 11815
rect 27445 11781 27479 11815
rect 29469 11781 29503 11815
rect 29669 11781 29703 11815
rect 35173 11781 35207 11815
rect 38117 11781 38151 11815
rect 1777 11713 1811 11747
rect 2421 11713 2455 11747
rect 5641 11713 5675 11747
rect 5733 11713 5767 11747
rect 6929 11713 6963 11747
rect 7297 11713 7331 11747
rect 8033 11713 8067 11747
rect 8217 11713 8251 11747
rect 8309 11713 8343 11747
rect 8401 11713 8435 11747
rect 9045 11713 9079 11747
rect 10057 11713 10091 11747
rect 10977 11713 11011 11747
rect 12265 11713 12299 11747
rect 12909 11713 12943 11747
rect 16129 11713 16163 11747
rect 17141 11713 17175 11747
rect 17289 11713 17323 11747
rect 17417 11713 17451 11747
rect 17647 11713 17681 11747
rect 18613 11713 18647 11747
rect 19441 11713 19475 11747
rect 21281 11713 21315 11747
rect 22017 11713 22051 11747
rect 22201 11713 22235 11747
rect 22385 11713 22419 11747
rect 23121 11713 23155 11747
rect 27169 11713 27203 11747
rect 30941 11713 30975 11747
rect 33885 11713 33919 11747
rect 38025 11713 38059 11747
rect 2697 11645 2731 11679
rect 5825 11645 5859 11679
rect 10149 11645 10183 11679
rect 10333 11645 10367 11679
rect 14933 11645 14967 11679
rect 15945 11645 15979 11679
rect 18705 11645 18739 11679
rect 18797 11645 18831 11679
rect 20637 11645 20671 11679
rect 23397 11645 23431 11679
rect 25789 11645 25823 11679
rect 25881 11645 25915 11679
rect 30481 11645 30515 11679
rect 31217 11645 31251 11679
rect 33149 11645 33183 11679
rect 33241 11645 33275 11679
rect 34897 11645 34931 11679
rect 4169 11577 4203 11611
rect 8585 11577 8619 11611
rect 9137 11577 9171 11611
rect 29837 11577 29871 11611
rect 30757 11577 30791 11611
rect 30849 11577 30883 11611
rect 1869 11509 1903 11543
rect 5273 11509 5307 11543
rect 6837 11509 6871 11543
rect 7021 11509 7055 11543
rect 9689 11509 9723 11543
rect 11069 11509 11103 11543
rect 12357 11509 12391 11543
rect 17785 11509 17819 11543
rect 18245 11509 18279 11543
rect 21373 11509 21407 11543
rect 22569 11509 22603 11543
rect 24869 11509 24903 11543
rect 29653 11509 29687 11543
rect 33977 11509 34011 11543
rect 2697 11305 2731 11339
rect 7941 11305 7975 11339
rect 8493 11305 8527 11339
rect 10885 11305 10919 11339
rect 16129 11305 16163 11339
rect 21741 11305 21775 11339
rect 23949 11305 23983 11339
rect 30757 11305 30791 11339
rect 34989 11305 35023 11339
rect 36277 11305 36311 11339
rect 6377 11237 6411 11271
rect 20177 11237 20211 11271
rect 27445 11237 27479 11271
rect 28733 11237 28767 11271
rect 29837 11237 29871 11271
rect 32045 11237 32079 11271
rect 34345 11237 34379 11271
rect 3157 11169 3191 11203
rect 3341 11169 3375 11203
rect 5733 11169 5767 11203
rect 9137 11169 9171 11203
rect 9413 11169 9447 11203
rect 11897 11169 11931 11203
rect 14381 11169 14415 11203
rect 14657 11169 14691 11203
rect 17325 11169 17359 11203
rect 18521 11169 18555 11203
rect 20729 11169 20763 11203
rect 22201 11169 22235 11203
rect 22385 11169 22419 11203
rect 25789 11169 25823 11203
rect 27905 11169 27939 11203
rect 27997 11169 28031 11203
rect 31217 11169 31251 11203
rect 31401 11169 31435 11203
rect 38577 11169 38611 11203
rect 2053 11101 2087 11135
rect 3985 11101 4019 11135
rect 6285 11101 6319 11135
rect 6929 11101 6963 11135
rect 7573 11101 7607 11135
rect 7757 11101 7791 11135
rect 8401 11101 8435 11135
rect 11713 11101 11747 11135
rect 13553 11101 13587 11135
rect 18245 11101 18279 11135
rect 19441 11101 19475 11135
rect 20545 11101 20579 11135
rect 23857 11101 23891 11135
rect 25513 11101 25547 11135
rect 26341 11101 26375 11135
rect 26525 11101 26559 11135
rect 26709 11101 26743 11135
rect 28641 11101 28675 11135
rect 29745 11101 29779 11135
rect 31953 11101 31987 11135
rect 32597 11101 32631 11135
rect 34897 11101 34931 11135
rect 35541 11101 35575 11135
rect 36185 11101 36219 11135
rect 36829 11101 36863 11135
rect 37565 11101 37599 11135
rect 1685 11033 1719 11067
rect 3065 11033 3099 11067
rect 4261 11033 4295 11067
rect 7021 11033 7055 11067
rect 13645 11033 13679 11067
rect 17233 11033 17267 11067
rect 20637 11033 20671 11067
rect 23029 11033 23063 11067
rect 23213 11033 23247 11067
rect 26617 11033 26651 11067
rect 27445 11033 27479 11067
rect 31125 11033 31159 11067
rect 32873 11033 32907 11067
rect 35633 11033 35667 11067
rect 37657 11033 37691 11067
rect 38301 11033 38335 11067
rect 16773 10965 16807 10999
rect 17141 10965 17175 10999
rect 19533 10965 19567 10999
rect 22109 10965 22143 10999
rect 25145 10965 25179 10999
rect 25605 10965 25639 10999
rect 26893 10965 26927 10999
rect 28181 10965 28215 10999
rect 36921 10965 36955 10999
rect 2145 10761 2179 10795
rect 5841 10761 5875 10795
rect 7037 10761 7071 10795
rect 14473 10761 14507 10795
rect 15393 10761 15427 10795
rect 17233 10761 17267 10795
rect 17325 10761 17359 10795
rect 19809 10761 19843 10795
rect 22109 10761 22143 10795
rect 25513 10761 25547 10795
rect 27169 10761 27203 10795
rect 30573 10761 30607 10795
rect 31033 10761 31067 10795
rect 2053 10693 2087 10727
rect 5641 10693 5675 10727
rect 6837 10693 6871 10727
rect 7941 10693 7975 10727
rect 9689 10693 9723 10727
rect 10425 10693 10459 10727
rect 13001 10693 13035 10727
rect 18337 10693 18371 10727
rect 25145 10693 25179 10727
rect 25345 10693 25379 10727
rect 29101 10693 29135 10727
rect 32597 10693 32631 10727
rect 2881 10625 2915 10659
rect 7665 10625 7699 10659
rect 10149 10625 10183 10659
rect 10333 10625 10367 10659
rect 10517 10625 10551 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 15485 10625 15519 10659
rect 20361 10625 20395 10659
rect 22017 10625 22051 10659
rect 25973 10625 26007 10659
rect 26066 10625 26100 10659
rect 26249 10625 26283 10659
rect 26341 10625 26375 10659
rect 26479 10625 26513 10659
rect 27537 10625 27571 10659
rect 27629 10625 27663 10659
rect 31401 10625 31435 10659
rect 34529 10625 34563 10659
rect 36737 10625 36771 10659
rect 37473 10625 37507 10659
rect 38117 10625 38151 10659
rect 3157 10557 3191 10591
rect 12725 10557 12759 10591
rect 15577 10557 15611 10591
rect 17417 10557 17451 10591
rect 18061 10557 18095 10591
rect 20913 10557 20947 10591
rect 22661 10557 22695 10591
rect 22937 10557 22971 10591
rect 24685 10557 24719 10591
rect 27721 10557 27755 10591
rect 28825 10557 28859 10591
rect 31493 10557 31527 10591
rect 31585 10557 31619 10591
rect 32321 10557 32355 10591
rect 34805 10557 34839 10591
rect 6009 10489 6043 10523
rect 16865 10489 16899 10523
rect 26617 10489 26651 10523
rect 4629 10421 4663 10455
rect 5825 10421 5859 10455
rect 7021 10421 7055 10455
rect 7205 10421 7239 10455
rect 10701 10421 10735 10455
rect 11713 10421 11747 10455
rect 12081 10421 12115 10455
rect 15025 10421 15059 10455
rect 25329 10421 25363 10455
rect 34069 10421 34103 10455
rect 36277 10421 36311 10455
rect 36829 10421 36863 10455
rect 37565 10421 37599 10455
rect 38209 10421 38243 10455
rect 5641 10217 5675 10251
rect 8585 10217 8619 10251
rect 12541 10217 12575 10251
rect 14381 10217 14415 10251
rect 15025 10217 15059 10251
rect 18521 10217 18555 10251
rect 26985 10217 27019 10251
rect 30389 10217 30423 10251
rect 31677 10217 31711 10251
rect 32965 10217 32999 10251
rect 38577 10217 38611 10251
rect 13001 10149 13035 10183
rect 25697 10149 25731 10183
rect 31953 10149 31987 10183
rect 4813 10081 4847 10115
rect 13461 10081 13495 10115
rect 13645 10081 13679 10115
rect 15577 10081 15611 10115
rect 17049 10081 17083 10115
rect 19809 10081 19843 10115
rect 20637 10081 20671 10115
rect 20913 10081 20947 10115
rect 23581 10081 23615 10115
rect 23673 10081 23707 10115
rect 31033 10081 31067 10115
rect 31677 10081 31711 10115
rect 34897 10081 34931 10115
rect 2329 10013 2363 10047
rect 3433 10013 3467 10047
rect 5549 10013 5583 10047
rect 6193 10013 6227 10047
rect 6837 10013 6871 10047
rect 9597 10013 9631 10047
rect 11989 10013 12023 10047
rect 12265 10013 12299 10047
rect 12357 10013 12391 10047
rect 13369 10013 13403 10047
rect 14289 10013 14323 10047
rect 16773 10013 16807 10047
rect 19533 10013 19567 10047
rect 22661 10013 22695 10047
rect 23489 10013 23523 10047
rect 24685 10013 24719 10047
rect 24797 10023 24831 10057
rect 26433 10013 26467 10047
rect 28549 10013 28583 10047
rect 28642 10013 28676 10047
rect 28917 10013 28951 10047
rect 29033 10013 29067 10047
rect 29745 10013 29779 10047
rect 30757 10013 30791 10047
rect 31585 10013 31619 10047
rect 32413 10013 32447 10047
rect 32781 10013 32815 10047
rect 33425 10013 33459 10047
rect 33793 10013 33827 10047
rect 37381 10013 37415 10047
rect 38393 10013 38427 10047
rect 1685 9945 1719 9979
rect 2237 9945 2271 9979
rect 2605 9945 2639 9979
rect 3249 9945 3283 9979
rect 4629 9945 4663 9979
rect 7113 9945 7147 9979
rect 9873 9945 9907 9979
rect 12173 9945 12207 9979
rect 15393 9945 15427 9979
rect 25697 9945 25731 9979
rect 26157 9945 26191 9979
rect 27261 9945 27295 9979
rect 27445 9945 27479 9979
rect 27537 9945 27571 9979
rect 28825 9945 28859 9979
rect 32597 9945 32631 9979
rect 32689 9945 32723 9979
rect 33609 9945 33643 9979
rect 33701 9945 33735 9979
rect 35173 9945 35207 9979
rect 36921 9945 36955 9979
rect 1777 9877 1811 9911
rect 4169 9877 4203 9911
rect 4537 9877 4571 9911
rect 6285 9877 6319 9911
rect 9321 9877 9355 9911
rect 11345 9877 11379 9911
rect 15485 9877 15519 9911
rect 23121 9877 23155 9911
rect 24961 9877 24995 9911
rect 26249 9877 26283 9911
rect 29193 9877 29227 9911
rect 29837 9877 29871 9911
rect 30849 9877 30883 9911
rect 33977 9877 34011 9911
rect 37473 9877 37507 9911
rect 13645 9673 13679 9707
rect 29285 9673 29319 9707
rect 29377 9673 29411 9707
rect 4905 9605 4939 9639
rect 5641 9605 5675 9639
rect 14105 9605 14139 9639
rect 15209 9605 15243 9639
rect 16221 9605 16255 9639
rect 17601 9605 17635 9639
rect 17785 9605 17819 9639
rect 17877 9605 17911 9639
rect 21189 9605 21223 9639
rect 22109 9605 22143 9639
rect 24041 9605 24075 9639
rect 27905 9605 27939 9639
rect 27997 9605 28031 9639
rect 28825 9605 28859 9639
rect 33517 9605 33551 9639
rect 36829 9605 36863 9639
rect 1593 9537 1627 9571
rect 4813 9537 4847 9571
rect 5457 9537 5491 9571
rect 5733 9537 5767 9571
rect 5825 9537 5859 9571
rect 11805 9537 11839 9571
rect 12541 9537 12575 9571
rect 14013 9537 14047 9571
rect 15301 9537 15335 9571
rect 16129 9537 16163 9571
rect 18705 9537 18739 9571
rect 20913 9537 20947 9571
rect 21097 9537 21131 9571
rect 21281 9537 21315 9571
rect 22256 9537 22290 9571
rect 23765 9537 23799 9571
rect 26065 9537 26099 9571
rect 26249 9537 26283 9571
rect 26341 9537 26375 9571
rect 26433 9537 26467 9571
rect 32321 9537 32355 9571
rect 35633 9537 35667 9571
rect 36185 9537 36219 9571
rect 36737 9537 36771 9571
rect 37473 9537 37507 9571
rect 38117 9537 38151 9571
rect 2421 9469 2455 9503
rect 2697 9469 2731 9503
rect 7113 9469 7147 9503
rect 7389 9469 7423 9503
rect 9321 9469 9355 9503
rect 9597 9469 9631 9503
rect 13093 9469 13127 9503
rect 14289 9469 14323 9503
rect 15393 9469 15427 9503
rect 18981 9469 19015 9503
rect 22477 9469 22511 9503
rect 22753 9469 22787 9503
rect 28181 9469 28215 9503
rect 29561 9469 29595 9503
rect 30021 9469 30055 9503
rect 30297 9469 30331 9503
rect 31769 9469 31803 9503
rect 32597 9469 32631 9503
rect 33241 9469 33275 9503
rect 11069 9401 11103 9435
rect 14841 9401 14875 9435
rect 21465 9401 21499 9435
rect 26617 9401 26651 9435
rect 28825 9401 28859 9435
rect 37565 9401 37599 9435
rect 1777 9333 1811 9367
rect 4169 9333 4203 9367
rect 6009 9333 6043 9367
rect 8861 9333 8895 9367
rect 11897 9333 11931 9367
rect 17325 9333 17359 9367
rect 20453 9333 20487 9367
rect 22385 9333 22419 9367
rect 25513 9333 25547 9367
rect 27537 9333 27571 9367
rect 34989 9333 35023 9367
rect 38209 9333 38243 9367
rect 2329 9129 2363 9163
rect 4248 9129 4282 9163
rect 6561 9129 6595 9163
rect 8401 9129 8435 9163
rect 9413 9129 9447 9163
rect 12817 9129 12851 9163
rect 26341 9129 26375 9163
rect 34897 9129 34931 9163
rect 36185 9129 36219 9163
rect 38577 9129 38611 9163
rect 12357 9061 12391 9095
rect 22845 9061 22879 9095
rect 29009 9061 29043 9095
rect 30297 9061 30331 9095
rect 2881 8993 2915 9027
rect 3985 8993 4019 9027
rect 7113 8993 7147 9027
rect 10057 8993 10091 9027
rect 10609 8993 10643 9027
rect 13461 8993 13495 9027
rect 14950 8993 14984 9027
rect 15485 8993 15519 9027
rect 20545 8993 20579 9027
rect 23581 8993 23615 9027
rect 24593 8993 24627 9027
rect 27537 8993 27571 9027
rect 30757 8993 30791 9027
rect 35357 8993 35391 9027
rect 35541 8993 35575 9027
rect 36829 8993 36863 9027
rect 1593 8925 1627 8959
rect 2697 8925 2731 8959
rect 6929 8925 6963 8959
rect 7021 8925 7055 8959
rect 7757 8925 7791 8959
rect 7850 8925 7884 8959
rect 8125 8925 8159 8959
rect 8222 8925 8256 8959
rect 9781 8925 9815 8959
rect 13185 8925 13219 8959
rect 14381 8925 14415 8959
rect 14801 8925 14835 8959
rect 18337 8925 18371 8959
rect 18521 8925 18555 8959
rect 18705 8925 18739 8959
rect 19441 8925 19475 8959
rect 19534 8925 19568 8959
rect 19717 8925 19751 8959
rect 19947 8925 19981 8959
rect 23305 8925 23339 8959
rect 27261 8925 27295 8959
rect 29745 8925 29779 8959
rect 30113 8925 30147 8959
rect 33517 8925 33551 8959
rect 33701 8925 33735 8959
rect 33885 8925 33919 8959
rect 35265 8925 35299 8959
rect 36093 8925 36127 8959
rect 2789 8857 2823 8891
rect 8033 8857 8067 8891
rect 9873 8857 9907 8891
rect 10885 8857 10919 8891
rect 13277 8857 13311 8891
rect 14565 8857 14599 8891
rect 14657 8857 14691 8891
rect 15761 8857 15795 8891
rect 17509 8857 17543 8891
rect 18613 8857 18647 8891
rect 19809 8857 19843 8891
rect 20821 8857 20855 8891
rect 22845 8857 22879 8891
rect 24869 8857 24903 8891
rect 29929 8857 29963 8891
rect 30021 8857 30055 8891
rect 31033 8857 31067 8891
rect 33793 8857 33827 8891
rect 37105 8857 37139 8891
rect 1777 8789 1811 8823
rect 5733 8789 5767 8823
rect 18889 8789 18923 8823
rect 20085 8789 20119 8823
rect 22293 8789 22327 8823
rect 23397 8789 23431 8823
rect 32505 8789 32539 8823
rect 34069 8789 34103 8823
rect 2881 8585 2915 8619
rect 3249 8585 3283 8619
rect 14105 8585 14139 8619
rect 14565 8585 14599 8619
rect 20729 8585 20763 8619
rect 22017 8585 22051 8619
rect 22385 8585 22419 8619
rect 22477 8585 22511 8619
rect 23581 8585 23615 8619
rect 25789 8585 25823 8619
rect 26157 8585 26191 8619
rect 26249 8585 26283 8619
rect 28917 8585 28951 8619
rect 32321 8585 32355 8619
rect 32781 8585 32815 8619
rect 33977 8585 34011 8619
rect 37473 8585 37507 8619
rect 37933 8585 37967 8619
rect 4537 8517 4571 8551
rect 7021 8517 7055 8551
rect 8585 8517 8619 8551
rect 10333 8517 10367 8551
rect 10793 8517 10827 8551
rect 11009 8517 11043 8551
rect 13185 8517 13219 8551
rect 14473 8517 14507 8551
rect 17141 8517 17175 8551
rect 27445 8517 27479 8551
rect 31033 8517 31067 8551
rect 32689 8517 32723 8551
rect 1593 8449 1627 8483
rect 1869 8449 1903 8483
rect 3341 8449 3375 8483
rect 4261 8449 4295 8483
rect 6929 8449 6963 8483
rect 11897 8449 11931 8483
rect 12265 8449 12299 8483
rect 12449 8449 12483 8483
rect 12725 8449 12759 8483
rect 15945 8449 15979 8483
rect 16037 8449 16071 8483
rect 16865 8449 16899 8483
rect 18889 8449 18923 8483
rect 19717 8449 19751 8483
rect 21097 8449 21131 8483
rect 23305 8449 23339 8483
rect 24685 8449 24719 8483
rect 25237 8449 25271 8483
rect 29837 8449 29871 8483
rect 31125 8449 31159 8483
rect 33885 8449 33919 8483
rect 34897 8449 34931 8483
rect 36001 8449 36035 8483
rect 36185 8449 36219 8483
rect 37841 8449 37875 8483
rect 3433 8381 3467 8415
rect 6009 8381 6043 8415
rect 7113 8381 7147 8415
rect 8309 8381 8343 8415
rect 11713 8381 11747 8415
rect 14657 8381 14691 8415
rect 16221 8381 16255 8415
rect 19809 8381 19843 8415
rect 19993 8381 20027 8415
rect 21189 8381 21223 8415
rect 21373 8381 21407 8415
rect 22661 8381 22695 8415
rect 26433 8381 26467 8415
rect 27169 8381 27203 8415
rect 29929 8381 29963 8415
rect 30113 8381 30147 8415
rect 31217 8381 31251 8415
rect 32965 8381 32999 8415
rect 34069 8381 34103 8415
rect 35173 8381 35207 8415
rect 38025 8381 38059 8415
rect 6561 8313 6595 8347
rect 11161 8313 11195 8347
rect 15577 8313 15611 8347
rect 19349 8313 19383 8347
rect 29469 8313 29503 8347
rect 33517 8313 33551 8347
rect 36369 8313 36403 8347
rect 10977 8245 11011 8279
rect 30665 8245 30699 8279
rect 2145 8041 2179 8075
rect 3985 8041 4019 8075
rect 4445 8041 4479 8075
rect 13461 8041 13495 8075
rect 14381 8041 14415 8075
rect 17693 8041 17727 8075
rect 17877 8041 17911 8075
rect 18889 8041 18923 8075
rect 24593 8041 24627 8075
rect 30002 8041 30036 8075
rect 31493 8041 31527 8075
rect 33701 8041 33735 8075
rect 35081 8041 35115 8075
rect 2329 7973 2363 8007
rect 13645 7973 13679 8007
rect 37749 7973 37783 8007
rect 4077 7905 4111 7939
rect 5549 7905 5583 7939
rect 6285 7905 6319 7939
rect 9781 7905 9815 7939
rect 11069 7905 11103 7939
rect 12817 7905 12851 7939
rect 15669 7905 15703 7939
rect 16773 7905 16807 7939
rect 16865 7905 16899 7939
rect 23857 7905 23891 7939
rect 25237 7905 25271 7939
rect 27077 7905 27111 7939
rect 29745 7905 29779 7939
rect 31953 7905 31987 7939
rect 35173 7905 35207 7939
rect 36001 7905 36035 7939
rect 2789 7837 2823 7871
rect 3157 7837 3191 7871
rect 4261 7837 4295 7871
rect 5273 7837 5307 7871
rect 10793 7837 10827 7871
rect 14289 7837 14323 7871
rect 14933 7837 14967 7871
rect 18337 7837 18371 7871
rect 18705 7837 18739 7871
rect 19809 7837 19843 7871
rect 22109 7837 22143 7871
rect 25789 7837 25823 7871
rect 26157 7837 26191 7871
rect 26801 7837 26835 7871
rect 28825 7837 28859 7871
rect 34161 7837 34195 7871
rect 35081 7837 35115 7871
rect 35357 7837 35391 7871
rect 38485 7837 38519 7871
rect 1961 7769 1995 7803
rect 2177 7769 2211 7803
rect 2973 7769 3007 7803
rect 3065 7769 3099 7803
rect 3985 7769 4019 7803
rect 6561 7769 6595 7803
rect 9505 7769 9539 7803
rect 13277 7769 13311 7803
rect 16681 7769 16715 7803
rect 17509 7769 17543 7803
rect 18521 7769 18555 7803
rect 18613 7769 18647 7803
rect 20085 7769 20119 7803
rect 22477 7769 22511 7803
rect 23581 7769 23615 7803
rect 25053 7769 25087 7803
rect 25973 7769 26007 7803
rect 26065 7769 26099 7803
rect 32229 7769 32263 7803
rect 34253 7769 34287 7803
rect 36277 7769 36311 7803
rect 38669 7769 38703 7803
rect 3341 7701 3375 7735
rect 4905 7701 4939 7735
rect 5365 7701 5399 7735
rect 8033 7701 8067 7735
rect 9137 7701 9171 7735
rect 9597 7701 9631 7735
rect 13487 7701 13521 7735
rect 16313 7701 16347 7735
rect 17719 7701 17753 7735
rect 21557 7701 21591 7735
rect 23213 7701 23247 7735
rect 23673 7701 23707 7735
rect 24961 7701 24995 7735
rect 26341 7701 26375 7735
rect 35541 7701 35575 7735
rect 3341 7497 3375 7531
rect 5641 7497 5675 7531
rect 23397 7497 23431 7531
rect 23857 7497 23891 7531
rect 24895 7497 24929 7531
rect 27169 7497 27203 7531
rect 27629 7497 27663 7531
rect 30941 7497 30975 7531
rect 31309 7497 31343 7531
rect 34279 7497 34313 7531
rect 36921 7497 36955 7531
rect 37841 7497 37875 7531
rect 2973 7429 3007 7463
rect 9321 7429 9355 7463
rect 12081 7429 12115 7463
rect 12173 7429 12207 7463
rect 13093 7429 13127 7463
rect 14197 7429 14231 7463
rect 15945 7429 15979 7463
rect 18521 7429 18555 7463
rect 18737 7429 18771 7463
rect 22569 7429 22603 7463
rect 24685 7429 24719 7463
rect 25513 7429 25547 7463
rect 27537 7429 27571 7463
rect 34069 7429 34103 7463
rect 37933 7429 37967 7463
rect 2053 7361 2087 7395
rect 2789 7361 2823 7395
rect 3065 7361 3099 7395
rect 3157 7361 3191 7395
rect 4169 7361 4203 7395
rect 4353 7361 4387 7395
rect 4813 7361 4847 7395
rect 7113 7361 7147 7395
rect 10977 7361 11011 7395
rect 12909 7361 12943 7395
rect 13185 7361 13219 7395
rect 13277 7361 13311 7395
rect 13921 7361 13955 7395
rect 17693 7361 17727 7395
rect 17785 7361 17819 7395
rect 19349 7361 19383 7395
rect 22385 7361 22419 7395
rect 22661 7361 22695 7395
rect 22753 7361 22787 7395
rect 23765 7361 23799 7395
rect 28641 7361 28675 7395
rect 31401 7361 31435 7395
rect 32689 7361 32723 7395
rect 33517 7361 33551 7395
rect 35173 7361 35207 7395
rect 4077 7293 4111 7327
rect 5733 7293 5767 7327
rect 5825 7293 5859 7327
rect 7389 7293 7423 7327
rect 10057 7293 10091 7327
rect 12357 7293 12391 7327
rect 17877 7293 17911 7327
rect 19625 7293 19659 7327
rect 21373 7293 21407 7327
rect 24041 7293 24075 7327
rect 26249 7293 26283 7327
rect 27721 7293 27755 7327
rect 28917 7293 28951 7327
rect 30389 7293 30423 7327
rect 31585 7293 31619 7327
rect 35449 7293 35483 7327
rect 38025 7293 38059 7327
rect 11069 7225 11103 7259
rect 25053 7225 25087 7259
rect 34437 7225 34471 7259
rect 37473 7225 37507 7259
rect 2237 7157 2271 7191
rect 5273 7157 5307 7191
rect 8861 7157 8895 7191
rect 11713 7157 11747 7191
rect 13461 7157 13495 7191
rect 17325 7157 17359 7191
rect 18705 7157 18739 7191
rect 18889 7157 18923 7191
rect 22937 7157 22971 7191
rect 24869 7157 24903 7191
rect 34253 7157 34287 7191
rect 2053 6953 2087 6987
rect 5444 6953 5478 6987
rect 17030 6953 17064 6987
rect 21097 6953 21131 6987
rect 22280 6953 22314 6987
rect 28733 6953 28767 6987
rect 34161 6953 34195 6987
rect 37086 6953 37120 6987
rect 12817 6885 12851 6919
rect 3341 6817 3375 6851
rect 4629 6817 4663 6851
rect 5181 6817 5215 6851
rect 10517 6817 10551 6851
rect 11069 6817 11103 6851
rect 14381 6817 14415 6851
rect 16773 6817 16807 6851
rect 20453 6817 20487 6851
rect 22017 6817 22051 6851
rect 25145 6817 25179 6851
rect 27169 6817 27203 6851
rect 28917 6817 28951 6851
rect 30941 6817 30975 6851
rect 31125 6817 31159 6851
rect 35449 6817 35483 6851
rect 7665 6749 7699 6783
rect 9229 6749 9263 6783
rect 10241 6749 10275 6783
rect 13277 6749 13311 6783
rect 14289 6749 14323 6783
rect 14933 6749 14967 6783
rect 20269 6749 20303 6783
rect 21097 6749 21131 6783
rect 21189 6749 21223 6783
rect 27629 6749 27663 6783
rect 27777 6749 27811 6783
rect 27997 6749 28031 6783
rect 28094 6749 28128 6783
rect 29009 6749 29043 6783
rect 31677 6749 31711 6783
rect 31861 6749 31895 6783
rect 32045 6749 32079 6783
rect 32689 6749 32723 6783
rect 34069 6749 34103 6783
rect 35357 6749 35391 6783
rect 36093 6749 36127 6783
rect 36829 6749 36863 6783
rect 1869 6681 1903 6715
rect 2085 6681 2119 6715
rect 3065 6681 3099 6715
rect 8401 6681 8435 6715
rect 11345 6681 11379 6715
rect 13553 6681 13587 6715
rect 15669 6681 15703 6715
rect 18797 6681 18831 6715
rect 20361 6681 20395 6715
rect 24041 6681 24075 6715
rect 25421 6681 25455 6715
rect 27905 6681 27939 6715
rect 28733 6681 28767 6715
rect 29837 6681 29871 6715
rect 30849 6681 30883 6715
rect 31953 6681 31987 6715
rect 33517 6681 33551 6715
rect 36185 6681 36219 6715
rect 2237 6613 2271 6647
rect 2697 6613 2731 6647
rect 3157 6613 3191 6647
rect 3985 6613 4019 6647
rect 4353 6613 4387 6647
rect 4445 6613 4479 6647
rect 6929 6613 6963 6647
rect 9321 6613 9355 6647
rect 9873 6613 9907 6647
rect 10333 6613 10367 6647
rect 19901 6613 19935 6647
rect 21465 6613 21499 6647
rect 28273 6613 28307 6647
rect 29193 6613 29227 6647
rect 29929 6613 29963 6647
rect 30481 6613 30515 6647
rect 32229 6613 32263 6647
rect 34897 6613 34931 6647
rect 35265 6613 35299 6647
rect 38577 6613 38611 6647
rect 1777 6409 1811 6443
rect 5457 6409 5491 6443
rect 7113 6409 7147 6443
rect 12541 6409 12575 6443
rect 12633 6409 12667 6443
rect 13737 6409 13771 6443
rect 23397 6409 23431 6443
rect 23949 6409 23983 6443
rect 34161 6409 34195 6443
rect 36369 6409 36403 6443
rect 37473 6409 37507 6443
rect 37933 6409 37967 6443
rect 2697 6341 2731 6375
rect 3985 6341 4019 6375
rect 6745 6341 6779 6375
rect 9597 6341 9631 6375
rect 18521 6341 18555 6375
rect 20821 6341 20855 6375
rect 24317 6341 24351 6375
rect 24409 6341 24443 6375
rect 25513 6341 25547 6375
rect 27445 6341 27479 6375
rect 32689 6341 32723 6375
rect 33793 6341 33827 6375
rect 33885 6341 33919 6375
rect 1593 6273 1627 6307
rect 2789 6273 2823 6307
rect 6561 6273 6595 6307
rect 6837 6273 6871 6307
rect 6929 6273 6963 6307
rect 7562 6273 7596 6307
rect 10793 6273 10827 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 14565 6273 14599 6307
rect 17141 6273 17175 6307
rect 22109 6273 22143 6307
rect 23213 6273 23247 6307
rect 33655 6273 33689 6307
rect 33977 6273 34011 6307
rect 37841 6273 37875 6307
rect 2881 6205 2915 6239
rect 3709 6205 3743 6239
rect 7849 6205 7883 6239
rect 12817 6205 12851 6239
rect 13829 6205 13863 6239
rect 13921 6205 13955 6239
rect 14841 6205 14875 6239
rect 17417 6205 17451 6239
rect 18245 6205 18279 6239
rect 19993 6205 20027 6239
rect 20913 6205 20947 6239
rect 21097 6205 21131 6239
rect 22385 6205 22419 6239
rect 24593 6205 24627 6239
rect 26341 6205 26375 6239
rect 27169 6205 27203 6239
rect 29653 6205 29687 6239
rect 29929 6205 29963 6239
rect 32781 6205 32815 6239
rect 32965 6205 32999 6239
rect 34621 6205 34655 6239
rect 34897 6205 34931 6239
rect 38025 6205 38059 6239
rect 12173 6137 12207 6171
rect 16313 6137 16347 6171
rect 20453 6137 20487 6171
rect 32321 6137 32355 6171
rect 2329 6069 2363 6103
rect 10425 6069 10459 6103
rect 10701 6069 10735 6103
rect 10885 6069 10919 6103
rect 13369 6069 13403 6103
rect 28917 6069 28951 6103
rect 31401 6069 31435 6103
rect 7094 5865 7128 5899
rect 8585 5865 8619 5899
rect 10885 5865 10919 5899
rect 14473 5865 14507 5899
rect 19441 5865 19475 5899
rect 23213 5865 23247 5899
rect 23857 5865 23891 5899
rect 25145 5865 25179 5899
rect 26893 5865 26927 5899
rect 30941 5865 30975 5899
rect 38485 5865 38519 5899
rect 18153 5797 18187 5831
rect 19809 5797 19843 5831
rect 24041 5797 24075 5831
rect 26525 5797 26559 5831
rect 27721 5797 27755 5831
rect 1961 5729 1995 5763
rect 4629 5729 4663 5763
rect 9137 5729 9171 5763
rect 9413 5729 9447 5763
rect 12265 5729 12299 5763
rect 14933 5729 14967 5763
rect 15025 5729 15059 5763
rect 15945 5729 15979 5763
rect 17417 5729 17451 5763
rect 18705 5729 18739 5763
rect 20913 5729 20947 5763
rect 21465 5729 21499 5763
rect 25605 5729 25639 5763
rect 25789 5729 25823 5763
rect 26985 5729 27019 5763
rect 27077 5729 27111 5763
rect 28181 5729 28215 5763
rect 28365 5729 28399 5763
rect 30297 5729 30331 5763
rect 31493 5729 31527 5763
rect 32597 5729 32631 5763
rect 35909 5729 35943 5763
rect 37933 5729 37967 5763
rect 1685 5661 1719 5695
rect 3985 5661 4019 5695
rect 6837 5661 6871 5695
rect 11989 5661 12023 5695
rect 15669 5661 15703 5695
rect 18613 5661 18647 5695
rect 19441 5661 19475 5695
rect 19625 5661 19659 5695
rect 20637 5661 20671 5695
rect 20729 5661 20763 5695
rect 24869 5661 24903 5695
rect 25513 5661 25547 5695
rect 26801 5661 26835 5695
rect 27261 5661 27295 5695
rect 28089 5661 28123 5695
rect 31401 5661 31435 5695
rect 34897 5661 34931 5695
rect 35081 5661 35115 5695
rect 38393 5661 38427 5695
rect 4905 5593 4939 5627
rect 21741 5593 21775 5627
rect 23673 5593 23707 5627
rect 29009 5593 29043 5627
rect 32873 5593 32907 5627
rect 35265 5593 35299 5627
rect 36185 5593 36219 5627
rect 3433 5525 3467 5559
rect 4077 5525 4111 5559
rect 6377 5525 6411 5559
rect 13737 5525 13771 5559
rect 14841 5525 14875 5559
rect 18521 5525 18555 5559
rect 20269 5525 20303 5559
rect 23883 5525 23917 5559
rect 29101 5525 29135 5559
rect 29745 5525 29779 5559
rect 30113 5525 30147 5559
rect 30205 5525 30239 5559
rect 31309 5525 31343 5559
rect 34345 5525 34379 5559
rect 1777 5321 1811 5355
rect 8309 5321 8343 5355
rect 9689 5321 9723 5355
rect 10425 5321 10459 5355
rect 13461 5321 13495 5355
rect 14013 5321 14047 5355
rect 31677 5321 31711 5355
rect 35357 5321 35391 5355
rect 35817 5321 35851 5355
rect 36763 5321 36797 5355
rect 37565 5321 37599 5355
rect 4353 5253 4387 5287
rect 6009 5253 6043 5287
rect 17141 5253 17175 5287
rect 21373 5253 21407 5287
rect 22569 5253 22603 5287
rect 23765 5253 23799 5287
rect 27353 5253 27387 5287
rect 32597 5253 32631 5287
rect 36553 5253 36587 5287
rect 1593 5185 1627 5219
rect 5273 5185 5307 5219
rect 9597 5185 9631 5219
rect 10793 5185 10827 5219
rect 13921 5185 13955 5219
rect 16865 5185 16899 5219
rect 21281 5185 21315 5219
rect 22661 5185 22695 5219
rect 24869 5185 24903 5219
rect 27169 5185 27203 5219
rect 27445 5185 27479 5219
rect 27537 5185 27571 5219
rect 28181 5185 28215 5219
rect 30757 5185 30791 5219
rect 30849 5185 30883 5219
rect 31585 5185 31619 5219
rect 32413 5185 32447 5219
rect 33149 5185 33183 5219
rect 35725 5185 35759 5219
rect 37473 5185 37507 5219
rect 38117 5185 38151 5219
rect 2329 5117 2363 5151
rect 2605 5117 2639 5151
rect 5641 5117 5675 5151
rect 6561 5117 6595 5151
rect 6837 5117 6871 5151
rect 9781 5117 9815 5151
rect 10885 5117 10919 5151
rect 11069 5117 11103 5151
rect 11713 5117 11747 5151
rect 11989 5117 12023 5151
rect 14565 5117 14599 5151
rect 14841 5117 14875 5151
rect 18613 5117 18647 5151
rect 19073 5117 19107 5151
rect 19349 5117 19383 5151
rect 20821 5117 20855 5151
rect 22753 5117 22787 5151
rect 23857 5117 23891 5151
rect 23949 5117 23983 5151
rect 25145 5117 25179 5151
rect 26617 5117 26651 5151
rect 28457 5117 28491 5151
rect 30941 5117 30975 5151
rect 33425 5117 33459 5151
rect 34897 5117 34931 5151
rect 35909 5117 35943 5151
rect 38209 5117 38243 5151
rect 5549 5049 5583 5083
rect 9229 5049 9263 5083
rect 23397 5049 23431 5083
rect 36921 5049 36955 5083
rect 5411 4981 5445 5015
rect 16313 4981 16347 5015
rect 22201 4981 22235 5015
rect 27721 4981 27755 5015
rect 29929 4981 29963 5015
rect 30389 4981 30423 5015
rect 36737 4981 36771 5015
rect 4537 4777 4571 4811
rect 4997 4777 5031 4811
rect 7941 4777 7975 4811
rect 9597 4777 9631 4811
rect 11437 4777 11471 4811
rect 25789 4777 25823 4811
rect 26065 4777 26099 4811
rect 33793 4777 33827 4811
rect 36645 4777 36679 4811
rect 38577 4777 38611 4811
rect 10241 4709 10275 4743
rect 12817 4709 12851 4743
rect 18153 4709 18187 4743
rect 26157 4709 26191 4743
rect 26985 4709 27019 4743
rect 31493 4709 31527 4743
rect 37289 4709 37323 4743
rect 1869 4641 1903 4675
rect 3341 4641 3375 4675
rect 5457 4641 5491 4675
rect 5549 4641 5583 4675
rect 6193 4641 6227 4675
rect 8493 4641 8527 4675
rect 10885 4641 10919 4675
rect 11897 4641 11931 4675
rect 12081 4641 12115 4675
rect 13277 4641 13311 4675
rect 13461 4641 13495 4675
rect 15301 4641 15335 4675
rect 17049 4641 17083 4675
rect 18613 4641 18647 4675
rect 18797 4641 18831 4675
rect 19901 4641 19935 4675
rect 19993 4641 20027 4675
rect 20913 4641 20947 4675
rect 26249 4641 26283 4675
rect 27537 4641 27571 4675
rect 30021 4641 30055 4675
rect 32045 4641 32079 4675
rect 37933 4641 37967 4675
rect 1593 4573 1627 4607
rect 3985 4573 4019 4607
rect 4169 4573 4203 4607
rect 4261 4573 4295 4607
rect 4353 4573 4387 4607
rect 8401 4573 8435 4607
rect 9045 4573 9079 4607
rect 9413 4573 9447 4607
rect 9873 4573 9907 4607
rect 14289 4573 14323 4607
rect 14473 4573 14507 4607
rect 14657 4573 14691 4607
rect 20637 4573 20671 4607
rect 23213 4573 23247 4607
rect 23581 4573 23615 4607
rect 24685 4573 24719 4607
rect 26341 4573 26375 4607
rect 26525 4573 26559 4607
rect 27445 4573 27479 4607
rect 28181 4573 28215 4607
rect 28365 4573 28399 4607
rect 28549 4573 28583 4607
rect 29745 4573 29779 4607
rect 35449 4573 35483 4607
rect 36553 4573 36587 4607
rect 37197 4573 37231 4607
rect 37841 4573 37875 4607
rect 38485 4573 38519 4607
rect 6469 4505 6503 4539
rect 9229 4505 9263 4539
rect 9321 4505 9355 4539
rect 10701 4505 10735 4539
rect 14565 4505 14599 4539
rect 15577 4505 15611 4539
rect 22661 4505 22695 4539
rect 25237 4505 25271 4539
rect 27353 4505 27387 4539
rect 28457 4505 28491 4539
rect 32321 4505 32355 4539
rect 35817 4505 35851 4539
rect 5365 4437 5399 4471
rect 10609 4437 10643 4471
rect 11805 4437 11839 4471
rect 13185 4437 13219 4471
rect 14841 4437 14875 4471
rect 18521 4437 18555 4471
rect 19441 4437 19475 4471
rect 19809 4437 19843 4471
rect 28733 4437 28767 4471
rect 5641 4233 5675 4267
rect 8033 4233 8067 4267
rect 9229 4233 9263 4267
rect 24041 4233 24075 4267
rect 24961 4233 24995 4267
rect 26065 4233 26099 4267
rect 35357 4233 35391 4267
rect 36553 4233 36587 4267
rect 1685 4165 1719 4199
rect 10609 4165 10643 4199
rect 10701 4165 10735 4199
rect 21097 4165 21131 4199
rect 35449 4165 35483 4199
rect 36645 4165 36679 4199
rect 6653 4097 6687 4131
rect 6837 4097 6871 4131
rect 6929 4097 6963 4131
rect 7021 4097 7055 4131
rect 9321 4097 9355 4131
rect 11713 4097 11747 4131
rect 12357 4097 12391 4131
rect 12541 4097 12575 4131
rect 12909 4097 12943 4131
rect 13093 4097 13127 4131
rect 13277 4097 13311 4131
rect 14289 4097 14323 4131
rect 16313 4097 16347 4131
rect 16957 4097 16991 4131
rect 17141 4097 17175 4131
rect 17233 4097 17267 4131
rect 17325 4097 17359 4131
rect 17969 4097 18003 4131
rect 21189 4097 21223 4131
rect 24869 4097 24903 4131
rect 27353 4097 27387 4131
rect 28365 4097 28399 4131
rect 28457 4097 28491 4131
rect 32321 4097 32355 4131
rect 37473 4097 37507 4131
rect 38117 4097 38151 4131
rect 2789 4029 2823 4063
rect 3065 4029 3099 4063
rect 4537 4029 4571 4063
rect 5733 4029 5767 4063
rect 5917 4029 5951 4063
rect 8125 4029 8159 4063
rect 8217 4029 8251 4063
rect 9505 4029 9539 4063
rect 10609 4029 10643 4063
rect 14565 4029 14599 4063
rect 18245 4029 18279 4063
rect 21373 4029 21407 4063
rect 22293 4029 22327 4063
rect 22569 4029 22603 4063
rect 25145 4029 25179 4063
rect 26157 4029 26191 4063
rect 26249 4029 26283 4063
rect 27169 4029 27203 4063
rect 28641 4029 28675 4063
rect 29469 4029 29503 4063
rect 29745 4029 29779 4063
rect 32597 4029 32631 4063
rect 35541 4029 35575 4063
rect 36737 4029 36771 4063
rect 7205 3961 7239 3995
rect 19717 3961 19751 3995
rect 37565 3961 37599 3995
rect 1777 3893 1811 3927
rect 5273 3893 5307 3927
rect 7665 3893 7699 3927
rect 8861 3893 8895 3927
rect 10149 3893 10183 3927
rect 11805 3893 11839 3927
rect 13737 3893 13771 3927
rect 17509 3893 17543 3927
rect 20729 3893 20763 3927
rect 24501 3893 24535 3927
rect 25697 3893 25731 3927
rect 27537 3893 27571 3927
rect 27997 3893 28031 3927
rect 31217 3893 31251 3927
rect 34069 3893 34103 3927
rect 34989 3893 35023 3927
rect 36185 3893 36219 3927
rect 38209 3893 38243 3927
rect 2697 3689 2731 3723
rect 3985 3689 4019 3723
rect 13645 3689 13679 3723
rect 16681 3689 16715 3723
rect 18889 3689 18923 3723
rect 22385 3689 22419 3723
rect 27261 3689 27295 3723
rect 27445 3689 27479 3723
rect 29929 3689 29963 3723
rect 30836 3689 30870 3723
rect 32965 3689 32999 3723
rect 5549 3621 5583 3655
rect 6653 3621 6687 3655
rect 21189 3621 21223 3655
rect 27997 3621 28031 3655
rect 30113 3621 30147 3655
rect 32321 3621 32355 3655
rect 36645 3621 36679 3655
rect 1869 3553 1903 3587
rect 3341 3553 3375 3587
rect 4537 3553 4571 3587
rect 6009 3553 6043 3587
rect 7297 3553 7331 3587
rect 8493 3553 8527 3587
rect 10057 3553 10091 3587
rect 14933 3553 14967 3587
rect 15209 3553 15243 3587
rect 17141 3553 17175 3587
rect 19441 3553 19475 3587
rect 19717 3553 19751 3587
rect 22937 3553 22971 3587
rect 23857 3553 23891 3587
rect 24777 3553 24811 3587
rect 25053 3553 25087 3587
rect 27169 3553 27203 3587
rect 28641 3553 28675 3587
rect 30573 3553 30607 3587
rect 33517 3553 33551 3587
rect 34897 3553 34931 3587
rect 1593 3485 1627 3519
rect 3065 3485 3099 3519
rect 3157 3485 3191 3519
rect 4353 3485 4387 3519
rect 7941 3485 7975 3519
rect 9873 3485 9907 3519
rect 11345 3485 11379 3519
rect 13553 3485 13587 3519
rect 14289 3485 14323 3519
rect 23581 3485 23615 3519
rect 27261 3485 27295 3519
rect 33333 3485 33367 3519
rect 34161 3485 34195 3519
rect 37197 3485 37231 3519
rect 38485 3485 38519 3519
rect 6101 3417 6135 3451
rect 11621 3417 11655 3451
rect 17417 3417 17451 3451
rect 21741 3417 21775 3451
rect 22753 3417 22787 3451
rect 26985 3417 27019 3451
rect 28457 3417 28491 3451
rect 29745 3417 29779 3451
rect 29961 3417 29995 3451
rect 35173 3417 35207 3451
rect 37013 3417 37047 3451
rect 38669 3417 38703 3451
rect 4445 3349 4479 3383
rect 6009 3349 6043 3383
rect 7021 3349 7055 3383
rect 7113 3349 7147 3383
rect 13093 3349 13127 3383
rect 14381 3349 14415 3383
rect 21833 3349 21867 3383
rect 22845 3349 22879 3383
rect 26525 3349 26559 3383
rect 28365 3349 28399 3383
rect 33425 3349 33459 3383
rect 34253 3349 34287 3383
rect 37289 3349 37323 3383
rect 4629 3145 4663 3179
rect 5733 3145 5767 3179
rect 6929 3145 6963 3179
rect 7389 3145 7423 3179
rect 10333 3145 10367 3179
rect 11805 3145 11839 3179
rect 12173 3145 12207 3179
rect 12265 3145 12299 3179
rect 15393 3145 15427 3179
rect 21097 3145 21131 3179
rect 25973 3145 26007 3179
rect 27629 3145 27663 3179
rect 1869 3077 1903 3111
rect 4261 3077 4295 3111
rect 8861 3077 8895 3111
rect 10977 3077 11011 3111
rect 18889 3077 18923 3111
rect 19625 3077 19659 3111
rect 22293 3077 22327 3111
rect 26525 3077 26559 3111
rect 32505 3077 32539 3111
rect 32597 3077 32631 3111
rect 33425 3077 33459 3111
rect 34253 3077 34287 3111
rect 34805 3077 34839 3111
rect 38485 3077 38519 3111
rect 1593 3009 1627 3043
rect 4077 3009 4111 3043
rect 4353 3009 4387 3043
rect 4445 3009 4479 3043
rect 5641 3009 5675 3043
rect 6561 3009 6595 3043
rect 6745 3009 6779 3043
rect 7757 3009 7791 3043
rect 13001 3009 13035 3043
rect 13645 3009 13679 3043
rect 15945 3009 15979 3043
rect 16865 3009 16899 3043
rect 19349 3009 19383 3043
rect 24225 3009 24259 3043
rect 26433 3009 26467 3043
rect 27537 3009 27571 3043
rect 31033 3009 31067 3043
rect 32321 3009 32355 3043
rect 32689 3009 32723 3043
rect 33977 3009 34011 3043
rect 35081 3009 35115 3043
rect 37473 3009 37507 3043
rect 3617 2941 3651 2975
rect 5917 2941 5951 2975
rect 7849 2941 7883 2975
rect 7941 2941 7975 2975
rect 8585 2941 8619 2975
rect 12449 2941 12483 2975
rect 13921 2941 13955 2975
rect 17141 2941 17175 2975
rect 22017 2941 22051 2975
rect 24501 2941 24535 2975
rect 27813 2941 27847 2975
rect 28641 2941 28675 2975
rect 28917 2941 28951 2975
rect 31585 2941 31619 2975
rect 35357 2941 35391 2975
rect 36829 2941 36863 2975
rect 11161 2873 11195 2907
rect 27169 2873 27203 2907
rect 32873 2873 32907 2907
rect 38669 2873 38703 2907
rect 5273 2805 5307 2839
rect 13093 2805 13127 2839
rect 16037 2805 16071 2839
rect 23765 2805 23799 2839
rect 30389 2805 30423 2839
rect 33517 2805 33551 2839
rect 37565 2805 37599 2839
rect 4997 2601 5031 2635
rect 6009 2601 6043 2635
rect 16037 2601 16071 2635
rect 18613 2601 18647 2635
rect 21189 2601 21223 2635
rect 22556 2601 22590 2635
rect 26341 2601 26375 2635
rect 28917 2601 28951 2635
rect 30849 2601 30883 2635
rect 34069 2601 34103 2635
rect 8309 2533 8343 2567
rect 11805 2533 11839 2567
rect 24041 2533 24075 2567
rect 34989 2533 35023 2567
rect 2329 2465 2363 2499
rect 6561 2465 6595 2499
rect 9873 2465 9907 2499
rect 12357 2465 12391 2499
rect 14289 2465 14323 2499
rect 16865 2465 16899 2499
rect 17141 2465 17175 2499
rect 19809 2465 19843 2499
rect 22293 2465 22327 2499
rect 24593 2465 24627 2499
rect 27169 2465 27203 2499
rect 30021 2465 30055 2499
rect 32321 2465 32355 2499
rect 36093 2465 36127 2499
rect 2053 2397 2087 2431
rect 2973 2397 3007 2431
rect 4445 2397 4479 2431
rect 4813 2397 4847 2431
rect 5457 2397 5491 2431
rect 5825 2397 5859 2431
rect 9597 2397 9631 2431
rect 10977 2397 11011 2431
rect 13093 2397 13127 2431
rect 19441 2397 19475 2431
rect 29745 2397 29779 2431
rect 31585 2397 31619 2431
rect 34897 2397 34931 2431
rect 35357 2397 35391 2431
rect 37565 2397 37599 2431
rect 3249 2329 3283 2363
rect 4629 2329 4663 2363
rect 4721 2329 4755 2363
rect 5641 2329 5675 2363
rect 5733 2329 5767 2363
rect 6837 2329 6871 2363
rect 12081 2329 12115 2363
rect 13461 2329 13495 2363
rect 14565 2329 14599 2363
rect 21097 2329 21131 2363
rect 24869 2329 24903 2363
rect 27445 2329 27479 2363
rect 30757 2329 30791 2363
rect 32597 2329 32631 2363
rect 35633 2329 35667 2363
rect 36553 2329 36587 2363
rect 38485 2329 38519 2363
rect 38669 2329 38703 2363
rect 11069 2261 11103 2295
rect 12265 2261 12299 2295
rect 31677 2261 31711 2295
rect 36645 2261 36679 2295
rect 37657 2261 37691 2295
<< metal1 >>
rect 16114 28228 16120 28280
rect 16172 28268 16178 28280
rect 17126 28268 17132 28280
rect 16172 28240 17132 28268
rect 16172 28228 16178 28240
rect 17126 28228 17132 28240
rect 17184 28228 17190 28280
rect 2314 26800 2320 26852
rect 2372 26840 2378 26852
rect 23750 26840 23756 26852
rect 2372 26812 23756 26840
rect 2372 26800 2378 26812
rect 23750 26800 23756 26812
rect 23808 26800 23814 26852
rect 26878 26732 26884 26784
rect 26936 26772 26942 26784
rect 34146 26772 34152 26784
rect 26936 26744 34152 26772
rect 26936 26732 26942 26744
rect 34146 26732 34152 26744
rect 34204 26732 34210 26784
rect 1104 26682 39192 26704
rect 1104 26630 5711 26682
rect 5763 26630 5775 26682
rect 5827 26630 5839 26682
rect 5891 26630 5903 26682
rect 5955 26630 5967 26682
rect 6019 26630 15233 26682
rect 15285 26630 15297 26682
rect 15349 26630 15361 26682
rect 15413 26630 15425 26682
rect 15477 26630 15489 26682
rect 15541 26630 24755 26682
rect 24807 26630 24819 26682
rect 24871 26630 24883 26682
rect 24935 26630 24947 26682
rect 24999 26630 25011 26682
rect 25063 26630 34277 26682
rect 34329 26630 34341 26682
rect 34393 26630 34405 26682
rect 34457 26630 34469 26682
rect 34521 26630 34533 26682
rect 34585 26630 39192 26682
rect 1104 26608 39192 26630
rect 658 26528 664 26580
rect 716 26568 722 26580
rect 3145 26571 3203 26577
rect 3145 26568 3157 26571
rect 716 26540 3157 26568
rect 716 26528 722 26540
rect 3145 26537 3157 26540
rect 3191 26537 3203 26571
rect 3145 26531 3203 26537
rect 8018 26528 8024 26580
rect 8076 26528 8082 26580
rect 26878 26568 26884 26580
rect 12406 26540 26884 26568
rect 6917 26503 6975 26509
rect 6917 26469 6929 26503
rect 6963 26500 6975 26503
rect 12406 26500 12434 26540
rect 26878 26528 26884 26540
rect 26936 26528 26942 26580
rect 27338 26528 27344 26580
rect 27396 26528 27402 26580
rect 27430 26528 27436 26580
rect 27488 26568 27494 26580
rect 29917 26571 29975 26577
rect 29917 26568 29929 26571
rect 27488 26540 29929 26568
rect 27488 26528 27494 26540
rect 29917 26537 29929 26540
rect 29963 26537 29975 26571
rect 29917 26531 29975 26537
rect 32490 26528 32496 26580
rect 32548 26528 32554 26580
rect 33594 26528 33600 26580
rect 33652 26568 33658 26580
rect 35069 26571 35127 26577
rect 35069 26568 35081 26571
rect 33652 26540 35081 26568
rect 33652 26528 33658 26540
rect 35069 26537 35081 26540
rect 35115 26537 35127 26571
rect 35069 26531 35127 26537
rect 37642 26528 37648 26580
rect 37700 26528 37706 26580
rect 6963 26472 12434 26500
rect 6963 26469 6975 26472
rect 6917 26463 6975 26469
rect 15562 26460 15568 26512
rect 15620 26500 15626 26512
rect 15620 26472 16068 26500
rect 15620 26460 15626 26472
rect 2314 26392 2320 26444
rect 2372 26392 2378 26444
rect 4249 26435 4307 26441
rect 4249 26401 4261 26435
rect 4295 26432 4307 26435
rect 13078 26432 13084 26444
rect 4295 26404 13084 26432
rect 4295 26401 4307 26404
rect 4249 26395 4307 26401
rect 13078 26392 13084 26404
rect 13136 26392 13142 26444
rect 13265 26435 13323 26441
rect 13265 26401 13277 26435
rect 13311 26432 13323 26435
rect 16040 26432 16068 26472
rect 16114 26460 16120 26512
rect 16172 26500 16178 26512
rect 16172 26472 20208 26500
rect 16172 26460 16178 26472
rect 18325 26435 18383 26441
rect 18325 26432 18337 26435
rect 13311 26404 15976 26432
rect 16040 26404 18337 26432
rect 13311 26401 13323 26404
rect 13265 26395 13323 26401
rect 2038 26324 2044 26376
rect 2096 26324 2102 26376
rect 3970 26324 3976 26376
rect 4028 26324 4034 26376
rect 6086 26324 6092 26376
rect 6144 26364 6150 26376
rect 6641 26367 6699 26373
rect 6641 26364 6653 26367
rect 6144 26336 6653 26364
rect 6144 26324 6150 26336
rect 6641 26333 6653 26336
rect 6687 26333 6699 26367
rect 6641 26327 6699 26333
rect 9122 26324 9128 26376
rect 9180 26324 9186 26376
rect 11330 26324 11336 26376
rect 11388 26364 11394 26376
rect 11701 26367 11759 26373
rect 11701 26364 11713 26367
rect 11388 26336 11713 26364
rect 11388 26324 11394 26336
rect 11701 26333 11713 26336
rect 11747 26333 11759 26367
rect 11701 26327 11759 26333
rect 12986 26324 12992 26376
rect 13044 26324 13050 26376
rect 14918 26324 14924 26376
rect 14976 26324 14982 26376
rect 15948 26364 15976 26404
rect 18325 26401 18337 26404
rect 18371 26401 18383 26435
rect 18325 26395 18383 26401
rect 16666 26364 16672 26376
rect 15948 26336 16672 26364
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 17126 26324 17132 26376
rect 17184 26324 17190 26376
rect 18138 26324 18144 26376
rect 18196 26324 18202 26376
rect 20180 26373 20208 26472
rect 20346 26460 20352 26512
rect 20404 26460 20410 26512
rect 34698 26500 34704 26512
rect 22066 26472 27292 26500
rect 20622 26392 20628 26444
rect 20680 26432 20686 26444
rect 22066 26432 22094 26472
rect 25593 26435 25651 26441
rect 25593 26432 25605 26435
rect 20680 26404 22094 26432
rect 23492 26404 25605 26432
rect 20680 26392 20686 26404
rect 20165 26367 20223 26373
rect 20165 26333 20177 26367
rect 20211 26333 20223 26367
rect 20165 26327 20223 26333
rect 22002 26324 22008 26376
rect 22060 26324 22066 26376
rect 23290 26324 23296 26376
rect 23348 26324 23354 26376
rect 3050 26256 3056 26308
rect 3108 26256 3114 26308
rect 7926 26256 7932 26308
rect 7984 26256 7990 26308
rect 9398 26256 9404 26308
rect 9456 26256 9462 26308
rect 15197 26299 15255 26305
rect 15197 26296 15209 26299
rect 14936 26268 15209 26296
rect 14936 26240 14964 26268
rect 15197 26265 15209 26268
rect 15243 26265 15255 26299
rect 15197 26259 15255 26265
rect 16942 26256 16948 26308
rect 17000 26256 17006 26308
rect 18506 26256 18512 26308
rect 18564 26296 18570 26308
rect 23492 26296 23520 26404
rect 25593 26401 25605 26404
rect 25639 26401 25651 26435
rect 25593 26395 25651 26401
rect 25130 26324 25136 26376
rect 25188 26364 25194 26376
rect 27264 26373 27292 26472
rect 27356 26472 34704 26500
rect 25317 26367 25375 26373
rect 25317 26364 25329 26367
rect 25188 26336 25329 26364
rect 25188 26324 25194 26336
rect 25317 26333 25329 26336
rect 25363 26333 25375 26367
rect 25317 26327 25375 26333
rect 27249 26367 27307 26373
rect 27249 26333 27261 26367
rect 27295 26333 27307 26367
rect 27249 26327 27307 26333
rect 18564 26268 23520 26296
rect 18564 26256 18570 26268
rect 23566 26256 23572 26308
rect 23624 26256 23630 26308
rect 27356 26296 27384 26472
rect 34698 26460 34704 26472
rect 34756 26460 34762 26512
rect 35526 26460 35532 26512
rect 35584 26500 35590 26512
rect 38473 26503 38531 26509
rect 38473 26500 38485 26503
rect 35584 26472 38485 26500
rect 35584 26460 35590 26472
rect 38473 26469 38485 26472
rect 38519 26469 38531 26503
rect 38473 26463 38531 26469
rect 27890 26392 27896 26444
rect 27948 26432 27954 26444
rect 27948 26404 28764 26432
rect 27948 26392 27954 26404
rect 28626 26373 28632 26376
rect 28445 26367 28503 26373
rect 28445 26333 28457 26367
rect 28491 26364 28503 26367
rect 28583 26367 28632 26373
rect 28491 26336 28525 26364
rect 28491 26333 28503 26336
rect 28445 26327 28503 26333
rect 28583 26333 28595 26367
rect 28629 26333 28632 26367
rect 28583 26327 28632 26333
rect 23676 26268 27384 26296
rect 11882 26188 11888 26240
rect 11940 26188 11946 26240
rect 14918 26188 14924 26240
rect 14976 26188 14982 26240
rect 22189 26231 22247 26237
rect 22189 26197 22201 26231
rect 22235 26228 22247 26231
rect 23676 26228 23704 26268
rect 28258 26256 28264 26308
rect 28316 26296 28322 26308
rect 28460 26296 28488 26327
rect 28626 26324 28632 26327
rect 28684 26324 28690 26376
rect 28736 26373 28764 26404
rect 29178 26392 29184 26444
rect 29236 26392 29242 26444
rect 36541 26435 36599 26441
rect 36541 26432 36553 26435
rect 29932 26404 36553 26432
rect 28721 26367 28779 26373
rect 28721 26333 28733 26367
rect 28767 26333 28779 26367
rect 28721 26327 28779 26333
rect 28994 26324 29000 26376
rect 29052 26364 29058 26376
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 29052 26336 29837 26364
rect 29052 26324 29058 26336
rect 29825 26333 29837 26336
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 29932 26296 29960 26404
rect 36541 26401 36553 26404
rect 36587 26401 36599 26435
rect 36541 26395 36599 26401
rect 30558 26324 30564 26376
rect 30616 26364 30622 26376
rect 30745 26367 30803 26373
rect 30745 26364 30757 26367
rect 30616 26336 30757 26364
rect 30616 26324 30622 26336
rect 30745 26333 30757 26336
rect 30791 26333 30803 26367
rect 30745 26327 30803 26333
rect 34606 26324 34612 26376
rect 34664 26364 34670 26376
rect 34977 26367 35035 26373
rect 34977 26364 34989 26367
rect 34664 26336 34989 26364
rect 34664 26324 34670 26336
rect 34977 26333 34989 26336
rect 35023 26333 35035 26367
rect 34977 26327 35035 26333
rect 36262 26324 36268 26376
rect 36320 26324 36326 26376
rect 38289 26367 38347 26373
rect 38289 26333 38301 26367
rect 38335 26364 38347 26367
rect 39390 26364 39396 26376
rect 38335 26336 39396 26364
rect 38335 26333 38347 26336
rect 38289 26327 38347 26333
rect 39390 26324 39396 26336
rect 39448 26324 39454 26376
rect 28316 26268 29960 26296
rect 28316 26256 28322 26268
rect 31110 26256 31116 26308
rect 31168 26256 31174 26308
rect 32398 26256 32404 26308
rect 32456 26256 32462 26308
rect 37550 26256 37556 26308
rect 37608 26296 37614 26308
rect 38013 26299 38071 26305
rect 38013 26296 38025 26299
rect 37608 26268 38025 26296
rect 37608 26256 37614 26268
rect 38013 26265 38025 26268
rect 38059 26265 38071 26299
rect 38013 26259 38071 26265
rect 22235 26200 23704 26228
rect 22235 26197 22247 26200
rect 22189 26191 22247 26197
rect 1104 26138 39352 26160
rect 1104 26086 10472 26138
rect 10524 26086 10536 26138
rect 10588 26086 10600 26138
rect 10652 26086 10664 26138
rect 10716 26086 10728 26138
rect 10780 26086 19994 26138
rect 20046 26086 20058 26138
rect 20110 26086 20122 26138
rect 20174 26086 20186 26138
rect 20238 26086 20250 26138
rect 20302 26086 29516 26138
rect 29568 26086 29580 26138
rect 29632 26086 29644 26138
rect 29696 26086 29708 26138
rect 29760 26086 29772 26138
rect 29824 26086 39038 26138
rect 39090 26086 39102 26138
rect 39154 26086 39166 26138
rect 39218 26086 39230 26138
rect 39282 26086 39294 26138
rect 39346 26086 39352 26138
rect 1104 26064 39352 26086
rect 934 25984 940 26036
rect 992 26024 998 26036
rect 1765 26027 1823 26033
rect 1765 26024 1777 26027
rect 992 25996 1777 26024
rect 992 25984 998 25996
rect 1765 25993 1777 25996
rect 1811 25993 1823 26027
rect 1765 25987 1823 25993
rect 18049 26027 18107 26033
rect 18049 25993 18061 26027
rect 18095 26024 18107 26027
rect 18874 26024 18880 26036
rect 18095 25996 18880 26024
rect 18095 25993 18107 25996
rect 18049 25987 18107 25993
rect 18874 25984 18880 25996
rect 18932 25984 18938 26036
rect 18138 25916 18144 25968
rect 18196 25956 18202 25968
rect 30190 25956 30196 25968
rect 18196 25928 30196 25956
rect 18196 25916 18202 25928
rect 30190 25916 30196 25928
rect 30248 25916 30254 25968
rect 38289 25959 38347 25965
rect 38289 25925 38301 25959
rect 38335 25956 38347 25959
rect 39482 25956 39488 25968
rect 38335 25928 39488 25956
rect 38335 25925 38347 25928
rect 38289 25919 38347 25925
rect 39482 25916 39488 25928
rect 39540 25916 39546 25968
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25888 1731 25891
rect 2130 25888 2136 25900
rect 1719 25860 2136 25888
rect 1719 25857 1731 25860
rect 1673 25851 1731 25857
rect 2130 25848 2136 25860
rect 2188 25848 2194 25900
rect 12986 25848 12992 25900
rect 13044 25888 13050 25900
rect 13173 25891 13231 25897
rect 13173 25888 13185 25891
rect 13044 25860 13185 25888
rect 13044 25848 13050 25860
rect 13173 25857 13185 25860
rect 13219 25888 13231 25891
rect 16117 25891 16175 25897
rect 16117 25888 16129 25891
rect 13219 25860 16129 25888
rect 13219 25857 13231 25860
rect 13173 25851 13231 25857
rect 16117 25857 16129 25860
rect 16163 25888 16175 25891
rect 16853 25891 16911 25897
rect 16853 25888 16865 25891
rect 16163 25860 16865 25888
rect 16163 25857 16175 25860
rect 16117 25851 16175 25857
rect 16853 25857 16865 25860
rect 16899 25857 16911 25891
rect 16853 25851 16911 25857
rect 17957 25891 18015 25897
rect 17957 25857 17969 25891
rect 18003 25888 18015 25891
rect 18506 25888 18512 25900
rect 18003 25860 18512 25888
rect 18003 25857 18015 25860
rect 17957 25851 18015 25857
rect 18506 25848 18512 25860
rect 18564 25848 18570 25900
rect 29365 25891 29423 25897
rect 29365 25857 29377 25891
rect 29411 25888 29423 25891
rect 30282 25888 30288 25900
rect 29411 25860 30288 25888
rect 29411 25857 29423 25860
rect 29365 25851 29423 25857
rect 30282 25848 30288 25860
rect 30340 25848 30346 25900
rect 37550 25848 37556 25900
rect 37608 25848 37614 25900
rect 8386 25780 8392 25832
rect 8444 25820 8450 25832
rect 9214 25820 9220 25832
rect 8444 25792 9220 25820
rect 8444 25780 8450 25792
rect 9214 25780 9220 25792
rect 9272 25820 9278 25832
rect 18230 25820 18236 25832
rect 9272 25792 18236 25820
rect 9272 25780 9278 25792
rect 18230 25780 18236 25792
rect 18288 25780 18294 25832
rect 14826 25712 14832 25764
rect 14884 25752 14890 25764
rect 34882 25752 34888 25764
rect 14884 25724 18000 25752
rect 14884 25712 14890 25724
rect 13265 25687 13323 25693
rect 13265 25653 13277 25687
rect 13311 25684 13323 25687
rect 13814 25684 13820 25696
rect 13311 25656 13820 25684
rect 13311 25653 13323 25656
rect 13265 25647 13323 25653
rect 13814 25644 13820 25656
rect 13872 25644 13878 25696
rect 16209 25687 16267 25693
rect 16209 25653 16221 25687
rect 16255 25684 16267 25687
rect 16758 25684 16764 25696
rect 16255 25656 16764 25684
rect 16255 25653 16267 25656
rect 16209 25647 16267 25653
rect 16758 25644 16764 25656
rect 16816 25644 16822 25696
rect 17034 25644 17040 25696
rect 17092 25644 17098 25696
rect 17126 25644 17132 25696
rect 17184 25684 17190 25696
rect 17589 25687 17647 25693
rect 17589 25684 17601 25687
rect 17184 25656 17601 25684
rect 17184 25644 17190 25656
rect 17589 25653 17601 25656
rect 17635 25653 17647 25687
rect 17972 25684 18000 25724
rect 22066 25724 34888 25752
rect 22066 25684 22094 25724
rect 34882 25712 34888 25724
rect 34940 25712 34946 25764
rect 17972 25656 22094 25684
rect 29365 25687 29423 25693
rect 17589 25647 17647 25653
rect 29365 25653 29377 25687
rect 29411 25684 29423 25687
rect 32766 25684 32772 25696
rect 29411 25656 32772 25684
rect 29411 25653 29423 25656
rect 29365 25647 29423 25653
rect 32766 25644 32772 25656
rect 32824 25644 32830 25696
rect 37642 25644 37648 25696
rect 37700 25644 37706 25696
rect 37918 25644 37924 25696
rect 37976 25684 37982 25696
rect 38381 25687 38439 25693
rect 38381 25684 38393 25687
rect 37976 25656 38393 25684
rect 37976 25644 37982 25656
rect 38381 25653 38393 25656
rect 38427 25653 38439 25687
rect 38381 25647 38439 25653
rect 1104 25594 39192 25616
rect 1104 25542 5711 25594
rect 5763 25542 5775 25594
rect 5827 25542 5839 25594
rect 5891 25542 5903 25594
rect 5955 25542 5967 25594
rect 6019 25542 15233 25594
rect 15285 25542 15297 25594
rect 15349 25542 15361 25594
rect 15413 25542 15425 25594
rect 15477 25542 15489 25594
rect 15541 25542 24755 25594
rect 24807 25542 24819 25594
rect 24871 25542 24883 25594
rect 24935 25542 24947 25594
rect 24999 25542 25011 25594
rect 25063 25542 34277 25594
rect 34329 25542 34341 25594
rect 34393 25542 34405 25594
rect 34457 25542 34469 25594
rect 34521 25542 34533 25594
rect 34585 25542 39192 25594
rect 1104 25520 39192 25542
rect 1026 25440 1032 25492
rect 1084 25480 1090 25492
rect 1765 25483 1823 25489
rect 1765 25480 1777 25483
rect 1084 25452 1777 25480
rect 1084 25440 1090 25452
rect 1765 25449 1777 25452
rect 1811 25449 1823 25483
rect 1765 25443 1823 25449
rect 8294 25440 8300 25492
rect 8352 25480 8358 25492
rect 8352 25452 18828 25480
rect 8352 25440 8358 25452
rect 7469 25347 7527 25353
rect 7469 25313 7481 25347
rect 7515 25344 7527 25347
rect 8386 25344 8392 25356
rect 7515 25316 8392 25344
rect 7515 25313 7527 25316
rect 7469 25307 7527 25313
rect 8386 25304 8392 25316
rect 8444 25304 8450 25356
rect 15657 25347 15715 25353
rect 15657 25313 15669 25347
rect 15703 25344 15715 25347
rect 17862 25344 17868 25356
rect 15703 25316 17868 25344
rect 15703 25313 15715 25316
rect 15657 25307 15715 25313
rect 17862 25304 17868 25316
rect 17920 25304 17926 25356
rect 18230 25304 18236 25356
rect 18288 25304 18294 25356
rect 1673 25279 1731 25285
rect 1673 25245 1685 25279
rect 1719 25276 1731 25279
rect 7926 25276 7932 25288
rect 1719 25248 7932 25276
rect 1719 25245 1731 25248
rect 1673 25239 1731 25245
rect 7926 25236 7932 25248
rect 7984 25236 7990 25288
rect 13906 25236 13912 25288
rect 13964 25276 13970 25288
rect 15381 25279 15439 25285
rect 15381 25276 15393 25279
rect 13964 25248 15393 25276
rect 13964 25236 13970 25248
rect 15381 25245 15393 25248
rect 15427 25245 15439 25279
rect 15381 25239 15439 25245
rect 18049 25279 18107 25285
rect 18049 25245 18061 25279
rect 18095 25276 18107 25279
rect 18138 25276 18144 25288
rect 18095 25248 18144 25276
rect 18095 25245 18107 25248
rect 18049 25239 18107 25245
rect 18138 25236 18144 25248
rect 18196 25236 18202 25288
rect 13081 25211 13139 25217
rect 13081 25177 13093 25211
rect 13127 25208 13139 25211
rect 14826 25208 14832 25220
rect 13127 25180 14832 25208
rect 13127 25177 13139 25180
rect 13081 25171 13139 25177
rect 14826 25168 14832 25180
rect 14884 25168 14890 25220
rect 18598 25208 18604 25220
rect 16882 25180 18604 25208
rect 18598 25168 18604 25180
rect 18656 25168 18662 25220
rect 6178 25100 6184 25152
rect 6236 25140 6242 25152
rect 6825 25143 6883 25149
rect 6825 25140 6837 25143
rect 6236 25112 6837 25140
rect 6236 25100 6242 25112
rect 6825 25109 6837 25112
rect 6871 25109 6883 25143
rect 6825 25103 6883 25109
rect 7190 25100 7196 25152
rect 7248 25100 7254 25152
rect 7285 25143 7343 25149
rect 7285 25109 7297 25143
rect 7331 25140 7343 25143
rect 7650 25140 7656 25152
rect 7331 25112 7656 25140
rect 7331 25109 7343 25112
rect 7285 25103 7343 25109
rect 7650 25100 7656 25112
rect 7708 25100 7714 25152
rect 13357 25143 13415 25149
rect 13357 25109 13369 25143
rect 13403 25140 13415 25143
rect 13538 25140 13544 25152
rect 13403 25112 13544 25140
rect 13403 25109 13415 25112
rect 13357 25103 13415 25109
rect 13538 25100 13544 25112
rect 13596 25100 13602 25152
rect 17129 25143 17187 25149
rect 17129 25109 17141 25143
rect 17175 25140 17187 25143
rect 18138 25140 18144 25152
rect 17175 25112 18144 25140
rect 17175 25109 17187 25112
rect 17129 25103 17187 25109
rect 18138 25100 18144 25112
rect 18196 25100 18202 25152
rect 18800 25140 18828 25452
rect 20898 25440 20904 25492
rect 20956 25480 20962 25492
rect 36633 25483 36691 25489
rect 20956 25452 35894 25480
rect 20956 25440 20962 25452
rect 29825 25415 29883 25421
rect 29825 25381 29837 25415
rect 29871 25412 29883 25415
rect 33318 25412 33324 25424
rect 29871 25384 33324 25412
rect 29871 25381 29883 25384
rect 29825 25375 29883 25381
rect 33318 25372 33324 25384
rect 33376 25372 33382 25424
rect 35866 25412 35894 25452
rect 36633 25449 36645 25483
rect 36679 25480 36691 25483
rect 36722 25480 36728 25492
rect 36679 25452 36728 25480
rect 36679 25449 36691 25452
rect 36633 25443 36691 25449
rect 36722 25440 36728 25452
rect 36780 25440 36786 25492
rect 38657 25415 38715 25421
rect 35866 25384 38516 25412
rect 27157 25347 27215 25353
rect 27157 25313 27169 25347
rect 27203 25344 27215 25347
rect 27798 25344 27804 25356
rect 27203 25316 27804 25344
rect 27203 25313 27215 25316
rect 27157 25307 27215 25313
rect 27798 25304 27804 25316
rect 27856 25304 27862 25356
rect 30190 25304 30196 25356
rect 30248 25344 30254 25356
rect 30377 25347 30435 25353
rect 30377 25344 30389 25347
rect 30248 25316 30389 25344
rect 30248 25304 30254 25316
rect 30377 25313 30389 25316
rect 30423 25313 30435 25347
rect 30377 25307 30435 25313
rect 25130 25236 25136 25288
rect 25188 25276 25194 25288
rect 26881 25279 26939 25285
rect 26881 25276 26893 25279
rect 25188 25248 26893 25276
rect 25188 25236 25194 25248
rect 26881 25245 26893 25248
rect 26927 25245 26939 25279
rect 26881 25239 26939 25245
rect 32677 25279 32735 25285
rect 32677 25245 32689 25279
rect 32723 25276 32735 25279
rect 36173 25279 36231 25285
rect 32723 25248 35894 25276
rect 32723 25245 32735 25248
rect 32677 25239 32735 25245
rect 30193 25211 30251 25217
rect 27264 25180 27646 25208
rect 27264 25140 27292 25180
rect 30193 25177 30205 25211
rect 30239 25208 30251 25211
rect 31110 25208 31116 25220
rect 30239 25180 31116 25208
rect 30239 25177 30251 25180
rect 30193 25171 30251 25177
rect 31110 25168 31116 25180
rect 31168 25168 31174 25220
rect 32582 25168 32588 25220
rect 32640 25208 32646 25220
rect 33045 25211 33103 25217
rect 33045 25208 33057 25211
rect 32640 25180 33057 25208
rect 32640 25168 32646 25180
rect 33045 25177 33057 25180
rect 33091 25177 33103 25211
rect 33045 25171 33103 25177
rect 18800 25112 27292 25140
rect 28442 25100 28448 25152
rect 28500 25140 28506 25152
rect 28629 25143 28687 25149
rect 28629 25140 28641 25143
rect 28500 25112 28641 25140
rect 28500 25100 28506 25112
rect 28629 25109 28641 25112
rect 28675 25109 28687 25143
rect 28629 25103 28687 25109
rect 28810 25100 28816 25152
rect 28868 25140 28874 25152
rect 30285 25143 30343 25149
rect 30285 25140 30297 25143
rect 28868 25112 30297 25140
rect 28868 25100 28874 25112
rect 30285 25109 30297 25112
rect 30331 25109 30343 25143
rect 35866 25140 35894 25248
rect 36173 25245 36185 25279
rect 36219 25276 36231 25279
rect 36262 25276 36268 25288
rect 36219 25248 36268 25276
rect 36219 25245 36231 25248
rect 36173 25239 36231 25245
rect 36262 25236 36268 25248
rect 36320 25236 36326 25288
rect 36446 25236 36452 25288
rect 36504 25276 36510 25288
rect 36541 25279 36599 25285
rect 36541 25276 36553 25279
rect 36504 25248 36553 25276
rect 36504 25236 36510 25248
rect 36541 25245 36553 25248
rect 36587 25245 36599 25279
rect 36541 25239 36599 25245
rect 36630 25236 36636 25288
rect 36688 25276 36694 25288
rect 38488 25285 38516 25384
rect 38657 25381 38669 25415
rect 38703 25412 38715 25415
rect 38930 25412 38936 25424
rect 38703 25384 38936 25412
rect 38703 25381 38715 25384
rect 38657 25375 38715 25381
rect 38930 25372 38936 25384
rect 38988 25372 38994 25424
rect 36725 25279 36783 25285
rect 36725 25276 36737 25279
rect 36688 25248 36737 25276
rect 36688 25236 36694 25248
rect 36725 25245 36737 25248
rect 36771 25245 36783 25279
rect 36725 25239 36783 25245
rect 38473 25279 38531 25285
rect 38473 25245 38485 25279
rect 38519 25245 38531 25279
rect 38473 25239 38531 25245
rect 36357 25143 36415 25149
rect 36357 25140 36369 25143
rect 35866 25112 36369 25140
rect 30285 25103 30343 25109
rect 36357 25109 36369 25112
rect 36403 25109 36415 25143
rect 36357 25103 36415 25109
rect 1104 25050 39352 25072
rect 1104 24998 10472 25050
rect 10524 24998 10536 25050
rect 10588 24998 10600 25050
rect 10652 24998 10664 25050
rect 10716 24998 10728 25050
rect 10780 24998 19994 25050
rect 20046 24998 20058 25050
rect 20110 24998 20122 25050
rect 20174 24998 20186 25050
rect 20238 24998 20250 25050
rect 20302 24998 29516 25050
rect 29568 24998 29580 25050
rect 29632 24998 29644 25050
rect 29696 24998 29708 25050
rect 29760 24998 29772 25050
rect 29824 24998 39038 25050
rect 39090 24998 39102 25050
rect 39154 24998 39166 25050
rect 39218 24998 39230 25050
rect 39282 24998 39294 25050
rect 39346 24998 39352 25050
rect 1104 24976 39352 24998
rect 18598 24896 18604 24948
rect 18656 24936 18662 24948
rect 28166 24936 28172 24948
rect 18656 24908 28172 24936
rect 18656 24896 18662 24908
rect 28166 24896 28172 24908
rect 28224 24896 28230 24948
rect 30374 24896 30380 24948
rect 30432 24936 30438 24948
rect 30432 24908 30604 24936
rect 30432 24896 30438 24908
rect 12989 24871 13047 24877
rect 12989 24837 13001 24871
rect 13035 24868 13047 24871
rect 14090 24868 14096 24880
rect 13035 24840 14096 24868
rect 13035 24837 13047 24840
rect 12989 24831 13047 24837
rect 14090 24828 14096 24840
rect 14148 24828 14154 24880
rect 17310 24828 17316 24880
rect 17368 24868 17374 24880
rect 17589 24871 17647 24877
rect 17589 24868 17601 24871
rect 17368 24840 17601 24868
rect 17368 24828 17374 24840
rect 17589 24837 17601 24840
rect 17635 24837 17647 24871
rect 17589 24831 17647 24837
rect 23569 24871 23627 24877
rect 23569 24837 23581 24871
rect 23615 24837 23627 24871
rect 30576 24868 30604 24908
rect 30926 24896 30932 24948
rect 30984 24936 30990 24948
rect 30984 24908 34836 24936
rect 30984 24896 30990 24908
rect 34808 24877 34836 24908
rect 34882 24896 34888 24948
rect 34940 24936 34946 24948
rect 34940 24908 36216 24936
rect 34940 24896 34946 24908
rect 36188 24877 36216 24908
rect 32585 24871 32643 24877
rect 32585 24868 32597 24871
rect 30576 24840 32597 24868
rect 23569 24831 23627 24837
rect 32585 24837 32597 24840
rect 32631 24837 32643 24871
rect 32585 24831 32643 24837
rect 34793 24871 34851 24877
rect 34793 24837 34805 24871
rect 34839 24837 34851 24871
rect 34793 24831 34851 24837
rect 36173 24871 36231 24877
rect 36173 24837 36185 24871
rect 36219 24837 36231 24871
rect 36173 24831 36231 24837
rect 12250 24760 12256 24812
rect 12308 24800 12314 24812
rect 14001 24803 14059 24809
rect 14001 24800 14013 24803
rect 12308 24772 14013 24800
rect 12308 24760 12314 24772
rect 14001 24769 14013 24772
rect 14047 24769 14059 24803
rect 14001 24763 14059 24769
rect 14826 24760 14832 24812
rect 14884 24760 14890 24812
rect 18138 24760 18144 24812
rect 18196 24760 18202 24812
rect 21634 24760 21640 24812
rect 21692 24800 21698 24812
rect 23584 24800 23612 24831
rect 36722 24828 36728 24880
rect 36780 24828 36786 24880
rect 25133 24803 25191 24809
rect 21692 24772 25084 24800
rect 21692 24760 21698 24772
rect 13078 24692 13084 24744
rect 13136 24692 13142 24744
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24732 13323 24735
rect 13538 24732 13544 24744
rect 13311 24704 13544 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 13538 24692 13544 24704
rect 13596 24692 13602 24744
rect 14734 24692 14740 24744
rect 14792 24732 14798 24744
rect 15013 24735 15071 24741
rect 15013 24732 15025 24735
rect 14792 24704 15025 24732
rect 14792 24692 14798 24704
rect 15013 24701 15025 24704
rect 15059 24701 15071 24735
rect 15013 24695 15071 24701
rect 17678 24692 17684 24744
rect 17736 24732 17742 24744
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 17736 24704 18061 24732
rect 17736 24692 17742 24704
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18049 24695 18107 24701
rect 23661 24735 23719 24741
rect 23661 24701 23673 24735
rect 23707 24732 23719 24735
rect 23750 24732 23756 24744
rect 23707 24704 23756 24732
rect 23707 24701 23719 24704
rect 23661 24695 23719 24701
rect 23750 24692 23756 24704
rect 23808 24692 23814 24744
rect 23842 24692 23848 24744
rect 23900 24692 23906 24744
rect 25056 24732 25084 24772
rect 25133 24769 25145 24803
rect 25179 24800 25191 24803
rect 25498 24800 25504 24812
rect 25179 24772 25504 24800
rect 25179 24769 25191 24772
rect 25133 24763 25191 24769
rect 25498 24760 25504 24772
rect 25556 24800 25562 24812
rect 28074 24800 28080 24812
rect 25556 24772 28080 24800
rect 25556 24760 25562 24772
rect 28074 24760 28080 24772
rect 28132 24760 28138 24812
rect 30282 24760 30288 24812
rect 30340 24800 30346 24812
rect 31018 24800 31024 24812
rect 30340 24772 31024 24800
rect 30340 24760 30346 24772
rect 31018 24760 31024 24772
rect 31076 24760 31082 24812
rect 25056 24704 31524 24732
rect 17402 24624 17408 24676
rect 17460 24664 17466 24676
rect 17589 24667 17647 24673
rect 17589 24664 17601 24667
rect 17460 24636 17601 24664
rect 17460 24624 17466 24636
rect 17589 24633 17601 24636
rect 17635 24633 17647 24667
rect 17589 24627 17647 24633
rect 24946 24624 24952 24676
rect 25004 24624 25010 24676
rect 30374 24664 30380 24676
rect 27448 24636 30380 24664
rect 12621 24599 12679 24605
rect 12621 24565 12633 24599
rect 12667 24596 12679 24599
rect 12710 24596 12716 24608
rect 12667 24568 12716 24596
rect 12667 24565 12679 24568
rect 12621 24559 12679 24565
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 14093 24599 14151 24605
rect 14093 24565 14105 24599
rect 14139 24596 14151 24599
rect 14182 24596 14188 24608
rect 14139 24568 14188 24596
rect 14139 24565 14151 24568
rect 14093 24559 14151 24565
rect 14182 24556 14188 24568
rect 14240 24556 14246 24608
rect 17034 24556 17040 24608
rect 17092 24596 17098 24608
rect 18325 24599 18383 24605
rect 18325 24596 18337 24599
rect 17092 24568 18337 24596
rect 17092 24556 17098 24568
rect 18325 24565 18337 24568
rect 18371 24565 18383 24599
rect 18325 24559 18383 24565
rect 23201 24599 23259 24605
rect 23201 24565 23213 24599
rect 23247 24596 23259 24599
rect 27448 24596 27476 24636
rect 30374 24624 30380 24636
rect 30432 24624 30438 24676
rect 23247 24568 27476 24596
rect 23247 24565 23259 24568
rect 23201 24559 23259 24565
rect 27614 24556 27620 24608
rect 27672 24596 27678 24608
rect 30101 24599 30159 24605
rect 30101 24596 30113 24599
rect 27672 24568 30113 24596
rect 27672 24556 27678 24568
rect 30101 24565 30113 24568
rect 30147 24565 30159 24599
rect 31496 24596 31524 24704
rect 31754 24692 31760 24744
rect 31812 24732 31818 24744
rect 32309 24735 32367 24741
rect 32309 24732 32321 24735
rect 31812 24704 32321 24732
rect 31812 24692 31818 24704
rect 32309 24701 32321 24704
rect 32355 24701 32367 24735
rect 32309 24695 32367 24701
rect 33704 24664 33732 24786
rect 34146 24760 34152 24812
rect 34204 24800 34210 24812
rect 35161 24803 35219 24809
rect 35161 24800 35173 24803
rect 34204 24772 35173 24800
rect 34204 24760 34210 24772
rect 35161 24769 35173 24772
rect 35207 24769 35219 24803
rect 35161 24763 35219 24769
rect 34698 24692 34704 24744
rect 34756 24692 34762 24744
rect 35176 24732 35204 24763
rect 35250 24760 35256 24812
rect 35308 24760 35314 24812
rect 35345 24803 35403 24809
rect 35345 24769 35357 24803
rect 35391 24800 35403 24803
rect 36262 24800 36268 24812
rect 35391 24772 36268 24800
rect 35391 24769 35403 24772
rect 35345 24763 35403 24769
rect 36262 24760 36268 24772
rect 36320 24800 36326 24812
rect 36538 24800 36544 24812
rect 36320 24772 36544 24800
rect 36320 24760 36326 24772
rect 36538 24760 36544 24772
rect 36596 24760 36602 24812
rect 36630 24760 36636 24812
rect 36688 24760 36694 24812
rect 38013 24803 38071 24809
rect 38013 24769 38025 24803
rect 38059 24800 38071 24803
rect 39390 24800 39396 24812
rect 38059 24772 39396 24800
rect 38059 24769 38071 24772
rect 38013 24763 38071 24769
rect 39390 24760 39396 24772
rect 39448 24760 39454 24812
rect 35894 24732 35900 24744
rect 35176 24704 35900 24732
rect 35894 24692 35900 24704
rect 35952 24692 35958 24744
rect 36078 24692 36084 24744
rect 36136 24732 36142 24744
rect 36446 24732 36452 24744
rect 36136 24704 36452 24732
rect 36136 24692 36142 24704
rect 36446 24692 36452 24704
rect 36504 24732 36510 24744
rect 36906 24732 36912 24744
rect 36504 24704 36912 24732
rect 36504 24692 36510 24704
rect 36906 24692 36912 24704
rect 36964 24692 36970 24744
rect 38286 24692 38292 24744
rect 38344 24692 38350 24744
rect 37642 24664 37648 24676
rect 33704 24636 37648 24664
rect 37642 24624 37648 24636
rect 37700 24624 37706 24676
rect 34057 24599 34115 24605
rect 34057 24596 34069 24599
rect 31496 24568 34069 24596
rect 30101 24559 30159 24565
rect 34057 24565 34069 24568
rect 34103 24565 34115 24599
rect 34057 24559 34115 24565
rect 35066 24556 35072 24608
rect 35124 24596 35130 24608
rect 36078 24596 36084 24608
rect 35124 24568 36084 24596
rect 35124 24556 35130 24568
rect 36078 24556 36084 24568
rect 36136 24556 36142 24608
rect 1104 24506 39192 24528
rect 1104 24454 5711 24506
rect 5763 24454 5775 24506
rect 5827 24454 5839 24506
rect 5891 24454 5903 24506
rect 5955 24454 5967 24506
rect 6019 24454 15233 24506
rect 15285 24454 15297 24506
rect 15349 24454 15361 24506
rect 15413 24454 15425 24506
rect 15477 24454 15489 24506
rect 15541 24454 24755 24506
rect 24807 24454 24819 24506
rect 24871 24454 24883 24506
rect 24935 24454 24947 24506
rect 24999 24454 25011 24506
rect 25063 24454 34277 24506
rect 34329 24454 34341 24506
rect 34393 24454 34405 24506
rect 34457 24454 34469 24506
rect 34521 24454 34533 24506
rect 34585 24454 39192 24506
rect 1104 24432 39192 24454
rect 8294 24352 8300 24404
rect 8352 24352 8358 24404
rect 12434 24352 12440 24404
rect 12492 24392 12498 24404
rect 15841 24395 15899 24401
rect 15841 24392 15853 24395
rect 12492 24364 15853 24392
rect 12492 24352 12498 24364
rect 15841 24361 15853 24364
rect 15887 24361 15899 24395
rect 15841 24355 15899 24361
rect 16209 24395 16267 24401
rect 16209 24361 16221 24395
rect 16255 24392 16267 24395
rect 16942 24392 16948 24404
rect 16255 24364 16948 24392
rect 16255 24361 16267 24364
rect 16209 24355 16267 24361
rect 16942 24352 16948 24364
rect 17000 24352 17006 24404
rect 17862 24352 17868 24404
rect 17920 24352 17926 24404
rect 28166 24352 28172 24404
rect 28224 24352 28230 24404
rect 34698 24352 34704 24404
rect 34756 24392 34762 24404
rect 35437 24395 35495 24401
rect 35437 24392 35449 24395
rect 34756 24364 35449 24392
rect 34756 24352 34762 24364
rect 35437 24361 35449 24364
rect 35483 24392 35495 24395
rect 36630 24392 36636 24404
rect 35483 24364 36636 24392
rect 35483 24361 35495 24364
rect 35437 24355 35495 24361
rect 36630 24352 36636 24364
rect 36688 24392 36694 24404
rect 36817 24395 36875 24401
rect 36817 24392 36829 24395
rect 36688 24364 36829 24392
rect 36688 24352 36694 24364
rect 36817 24361 36829 24364
rect 36863 24361 36875 24395
rect 36817 24355 36875 24361
rect 12621 24327 12679 24333
rect 12621 24293 12633 24327
rect 12667 24324 12679 24327
rect 12667 24296 14964 24324
rect 12667 24293 12679 24296
rect 12621 24287 12679 24293
rect 6178 24216 6184 24268
rect 6236 24216 6242 24268
rect 6546 24216 6552 24268
rect 6604 24256 6610 24268
rect 6604 24228 8248 24256
rect 6604 24216 6610 24228
rect 934 24148 940 24200
rect 992 24188 998 24200
rect 8220 24197 8248 24228
rect 11974 24216 11980 24268
rect 12032 24256 12038 24268
rect 13173 24259 13231 24265
rect 13173 24256 13185 24259
rect 12032 24228 13185 24256
rect 12032 24216 12038 24228
rect 13173 24225 13185 24228
rect 13219 24225 13231 24259
rect 13173 24219 13231 24225
rect 14734 24216 14740 24268
rect 14792 24256 14798 24268
rect 14829 24259 14887 24265
rect 14829 24256 14841 24259
rect 14792 24228 14841 24256
rect 14792 24216 14798 24228
rect 14829 24225 14841 24228
rect 14875 24225 14887 24259
rect 14936 24256 14964 24296
rect 15010 24284 15016 24336
rect 15068 24324 15074 24336
rect 19058 24324 19064 24336
rect 15068 24296 19064 24324
rect 15068 24284 15074 24296
rect 19058 24284 19064 24296
rect 19116 24284 19122 24336
rect 17218 24256 17224 24268
rect 14936 24228 17224 24256
rect 14829 24219 14887 24225
rect 17218 24216 17224 24228
rect 17276 24216 17282 24268
rect 18138 24216 18144 24268
rect 18196 24256 18202 24268
rect 18325 24259 18383 24265
rect 18325 24256 18337 24259
rect 18196 24228 18337 24256
rect 18196 24216 18202 24228
rect 18325 24225 18337 24228
rect 18371 24225 18383 24259
rect 18325 24219 18383 24225
rect 18509 24259 18567 24265
rect 18509 24225 18521 24259
rect 18555 24256 18567 24259
rect 18598 24256 18604 24268
rect 18555 24228 18604 24256
rect 18555 24225 18567 24228
rect 18509 24219 18567 24225
rect 18598 24216 18604 24228
rect 18656 24216 18662 24268
rect 20530 24216 20536 24268
rect 20588 24256 20594 24268
rect 26789 24259 26847 24265
rect 26789 24256 26801 24259
rect 20588 24228 26801 24256
rect 20588 24216 20594 24228
rect 26789 24225 26801 24228
rect 26835 24225 26847 24259
rect 26789 24219 26847 24225
rect 34974 24216 34980 24268
rect 35032 24256 35038 24268
rect 35529 24259 35587 24265
rect 35032 24228 35296 24256
rect 35032 24216 35038 24228
rect 1673 24191 1731 24197
rect 1673 24188 1685 24191
rect 992 24160 1685 24188
rect 992 24148 998 24160
rect 1673 24157 1685 24160
rect 1719 24157 1731 24191
rect 1673 24151 1731 24157
rect 5905 24191 5963 24197
rect 5905 24157 5917 24191
rect 5951 24157 5963 24191
rect 5905 24151 5963 24157
rect 8205 24191 8263 24197
rect 8205 24157 8217 24191
rect 8251 24157 8263 24191
rect 8205 24151 8263 24157
rect 2222 24080 2228 24132
rect 2280 24080 2286 24132
rect 5920 24120 5948 24151
rect 8478 24148 8484 24200
rect 8536 24188 8542 24200
rect 8536 24160 12434 24188
rect 8536 24148 8542 24160
rect 6086 24120 6092 24132
rect 5920 24092 6092 24120
rect 6086 24080 6092 24092
rect 6144 24080 6150 24132
rect 6638 24080 6644 24132
rect 6696 24080 6702 24132
rect 9309 24123 9367 24129
rect 9309 24089 9321 24123
rect 9355 24120 9367 24123
rect 10318 24120 10324 24132
rect 9355 24092 10324 24120
rect 9355 24089 9367 24092
rect 9309 24083 9367 24089
rect 10318 24080 10324 24092
rect 10376 24080 10382 24132
rect 12406 24120 12434 24160
rect 14918 24148 14924 24200
rect 14976 24188 14982 24200
rect 15194 24188 15200 24200
rect 14976 24160 15200 24188
rect 14976 24148 14982 24160
rect 15194 24148 15200 24160
rect 15252 24148 15258 24200
rect 15838 24148 15844 24200
rect 15896 24148 15902 24200
rect 16022 24148 16028 24200
rect 16080 24148 16086 24200
rect 26881 24191 26939 24197
rect 26881 24188 26893 24191
rect 19628 24160 26893 24188
rect 18233 24123 18291 24129
rect 18233 24120 18245 24123
rect 12406 24092 18245 24120
rect 18233 24089 18245 24092
rect 18279 24089 18291 24123
rect 18233 24083 18291 24089
rect 7650 24012 7656 24064
rect 7708 24012 7714 24064
rect 8938 24012 8944 24064
rect 8996 24052 9002 24064
rect 9401 24055 9459 24061
rect 9401 24052 9413 24055
rect 8996 24024 9413 24052
rect 8996 24012 9002 24024
rect 9401 24021 9413 24024
rect 9447 24021 9459 24055
rect 9401 24015 9459 24021
rect 12618 24012 12624 24064
rect 12676 24052 12682 24064
rect 12989 24055 13047 24061
rect 12989 24052 13001 24055
rect 12676 24024 13001 24052
rect 12676 24012 12682 24024
rect 12989 24021 13001 24024
rect 13035 24021 13047 24055
rect 12989 24015 13047 24021
rect 13081 24055 13139 24061
rect 13081 24021 13093 24055
rect 13127 24052 13139 24055
rect 13446 24052 13452 24064
rect 13127 24024 13452 24052
rect 13127 24021 13139 24024
rect 13081 24015 13139 24021
rect 13446 24012 13452 24024
rect 13504 24012 13510 24064
rect 14274 24012 14280 24064
rect 14332 24012 14338 24064
rect 14642 24012 14648 24064
rect 14700 24012 14706 24064
rect 14737 24055 14795 24061
rect 14737 24021 14749 24055
rect 14783 24052 14795 24055
rect 15102 24052 15108 24064
rect 14783 24024 15108 24052
rect 14783 24021 14795 24024
rect 14737 24015 14795 24021
rect 15102 24012 15108 24024
rect 15160 24012 15166 24064
rect 15194 24012 15200 24064
rect 15252 24052 15258 24064
rect 19628 24052 19656 24160
rect 26881 24157 26893 24160
rect 26927 24188 26939 24191
rect 26970 24188 26976 24200
rect 26927 24160 26976 24188
rect 26927 24157 26939 24160
rect 26881 24151 26939 24157
rect 26970 24148 26976 24160
rect 27028 24148 27034 24200
rect 27065 24191 27123 24197
rect 27065 24157 27077 24191
rect 27111 24188 27123 24191
rect 27706 24188 27712 24200
rect 27111 24160 27712 24188
rect 27111 24157 27123 24160
rect 27065 24151 27123 24157
rect 23842 24080 23848 24132
rect 23900 24120 23906 24132
rect 27080 24120 27108 24151
rect 27706 24148 27712 24160
rect 27764 24148 27770 24200
rect 28074 24148 28080 24200
rect 28132 24148 28138 24200
rect 28534 24148 28540 24200
rect 28592 24188 28598 24200
rect 31849 24191 31907 24197
rect 31849 24188 31861 24191
rect 28592 24160 31861 24188
rect 28592 24148 28598 24160
rect 31849 24157 31861 24160
rect 31895 24157 31907 24191
rect 31849 24151 31907 24157
rect 32582 24148 32588 24200
rect 32640 24148 32646 24200
rect 35066 24148 35072 24200
rect 35124 24148 35130 24200
rect 35268 24188 35296 24228
rect 35529 24225 35541 24259
rect 35575 24256 35587 24259
rect 35894 24256 35900 24268
rect 35575 24228 35900 24256
rect 35575 24225 35587 24228
rect 35529 24219 35587 24225
rect 35894 24216 35900 24228
rect 35952 24256 35958 24268
rect 35952 24228 36584 24256
rect 35952 24216 35958 24228
rect 36446 24188 36452 24200
rect 35268 24160 36452 24188
rect 36446 24148 36452 24160
rect 36504 24148 36510 24200
rect 36556 24197 36584 24228
rect 36541 24191 36599 24197
rect 36541 24157 36553 24191
rect 36587 24188 36599 24191
rect 36722 24188 36728 24200
rect 36587 24160 36728 24188
rect 36587 24157 36599 24160
rect 36541 24151 36599 24157
rect 36722 24148 36728 24160
rect 36780 24148 36786 24200
rect 36906 24148 36912 24200
rect 36964 24148 36970 24200
rect 23900 24092 27108 24120
rect 23900 24080 23906 24092
rect 27522 24080 27528 24132
rect 27580 24080 27586 24132
rect 32950 24080 32956 24132
rect 33008 24080 33014 24132
rect 15252 24024 19656 24052
rect 15252 24012 15258 24024
rect 19702 24012 19708 24064
rect 19760 24052 19766 24064
rect 27614 24052 27620 24064
rect 19760 24024 27620 24052
rect 19760 24012 19766 24024
rect 27614 24012 27620 24024
rect 27672 24012 27678 24064
rect 31941 24055 31999 24061
rect 31941 24021 31953 24055
rect 31987 24052 31999 24055
rect 32030 24052 32036 24064
rect 31987 24024 32036 24052
rect 31987 24021 31999 24024
rect 31941 24015 31999 24021
rect 32030 24012 32036 24024
rect 32088 24012 32094 24064
rect 35434 24012 35440 24064
rect 35492 24052 35498 24064
rect 35805 24055 35863 24061
rect 35805 24052 35817 24055
rect 35492 24024 35817 24052
rect 35492 24012 35498 24024
rect 35805 24021 35817 24024
rect 35851 24021 35863 24055
rect 35805 24015 35863 24021
rect 37090 24012 37096 24064
rect 37148 24012 37154 24064
rect 1104 23962 39352 23984
rect 1104 23910 10472 23962
rect 10524 23910 10536 23962
rect 10588 23910 10600 23962
rect 10652 23910 10664 23962
rect 10716 23910 10728 23962
rect 10780 23910 19994 23962
rect 20046 23910 20058 23962
rect 20110 23910 20122 23962
rect 20174 23910 20186 23962
rect 20238 23910 20250 23962
rect 20302 23910 29516 23962
rect 29568 23910 29580 23962
rect 29632 23910 29644 23962
rect 29696 23910 29708 23962
rect 29760 23910 29772 23962
rect 29824 23910 39038 23962
rect 39090 23910 39102 23962
rect 39154 23910 39166 23962
rect 39218 23910 39230 23962
rect 39282 23910 39294 23962
rect 39346 23910 39352 23962
rect 1104 23888 39352 23910
rect 5077 23851 5135 23857
rect 5077 23817 5089 23851
rect 5123 23848 5135 23851
rect 6638 23848 6644 23860
rect 5123 23820 6644 23848
rect 5123 23817 5135 23820
rect 5077 23811 5135 23817
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 7190 23808 7196 23860
rect 7248 23848 7254 23860
rect 7742 23848 7748 23860
rect 7248 23820 7748 23848
rect 7248 23808 7254 23820
rect 7742 23808 7748 23820
rect 7800 23848 7806 23860
rect 8205 23851 8263 23857
rect 8205 23848 8217 23851
rect 7800 23820 8217 23848
rect 7800 23808 7806 23820
rect 8205 23817 8217 23820
rect 8251 23817 8263 23851
rect 8205 23811 8263 23817
rect 12342 23808 12348 23860
rect 12400 23848 12406 23860
rect 13633 23851 13691 23857
rect 13633 23848 13645 23851
rect 12400 23820 13645 23848
rect 12400 23808 12406 23820
rect 13633 23817 13645 23820
rect 13679 23817 13691 23851
rect 13633 23811 13691 23817
rect 14093 23851 14151 23857
rect 14093 23817 14105 23851
rect 14139 23848 14151 23851
rect 15562 23848 15568 23860
rect 14139 23820 15568 23848
rect 14139 23817 14151 23820
rect 14093 23811 14151 23817
rect 15562 23808 15568 23820
rect 15620 23808 15626 23860
rect 30926 23848 30932 23860
rect 16546 23820 30932 23848
rect 11054 23780 11060 23792
rect 2746 23752 11060 23780
rect 2222 23536 2228 23588
rect 2280 23576 2286 23588
rect 2746 23576 2774 23752
rect 11054 23740 11060 23752
rect 11112 23740 11118 23792
rect 15010 23780 15016 23792
rect 12406 23752 15016 23780
rect 4154 23672 4160 23724
rect 4212 23712 4218 23724
rect 4985 23715 5043 23721
rect 4985 23712 4997 23715
rect 4212 23684 4997 23712
rect 4212 23672 4218 23684
rect 4985 23681 4997 23684
rect 5031 23681 5043 23715
rect 4985 23675 5043 23681
rect 6914 23672 6920 23724
rect 6972 23672 6978 23724
rect 7009 23715 7067 23721
rect 7009 23681 7021 23715
rect 7055 23712 7067 23715
rect 7834 23712 7840 23724
rect 7055 23684 7840 23712
rect 7055 23681 7067 23684
rect 7009 23675 7067 23681
rect 7834 23672 7840 23684
rect 7892 23672 7898 23724
rect 8110 23672 8116 23724
rect 8168 23712 8174 23724
rect 9125 23715 9183 23721
rect 8168 23684 8432 23712
rect 8168 23672 8174 23684
rect 4890 23604 4896 23656
rect 4948 23644 4954 23656
rect 7193 23647 7251 23653
rect 7193 23644 7205 23647
rect 4948 23616 7205 23644
rect 4948 23604 4954 23616
rect 7193 23613 7205 23616
rect 7239 23644 7251 23647
rect 7239 23616 8064 23644
rect 7239 23613 7251 23616
rect 7193 23607 7251 23613
rect 2280 23548 2774 23576
rect 8036 23576 8064 23616
rect 8202 23604 8208 23656
rect 8260 23644 8266 23656
rect 8404 23653 8432 23684
rect 9125 23681 9137 23715
rect 9171 23712 9183 23715
rect 12406 23712 12434 23752
rect 15010 23740 15016 23752
rect 15068 23740 15074 23792
rect 9171 23684 12434 23712
rect 9171 23681 9183 23684
rect 9125 23675 9183 23681
rect 12986 23672 12992 23724
rect 13044 23712 13050 23724
rect 13722 23712 13728 23724
rect 13044 23684 13728 23712
rect 13044 23672 13050 23684
rect 13722 23672 13728 23684
rect 13780 23672 13786 23724
rect 13998 23672 14004 23724
rect 14056 23672 14062 23724
rect 14829 23715 14887 23721
rect 14829 23681 14841 23715
rect 14875 23712 14887 23715
rect 16546 23712 16574 23820
rect 30926 23808 30932 23820
rect 30984 23848 30990 23860
rect 31294 23848 31300 23860
rect 30984 23820 31300 23848
rect 30984 23808 30990 23820
rect 31294 23808 31300 23820
rect 31352 23808 31358 23860
rect 25130 23780 25136 23792
rect 24872 23752 25136 23780
rect 14875 23684 16574 23712
rect 14875 23681 14887 23684
rect 14829 23675 14887 23681
rect 16850 23672 16856 23724
rect 16908 23712 16914 23724
rect 16945 23715 17003 23721
rect 16945 23712 16957 23715
rect 16908 23684 16957 23712
rect 16908 23672 16914 23684
rect 16945 23681 16957 23684
rect 16991 23712 17003 23715
rect 17310 23712 17316 23724
rect 16991 23684 17316 23712
rect 16991 23681 17003 23684
rect 16945 23675 17003 23681
rect 17310 23672 17316 23684
rect 17368 23672 17374 23724
rect 17402 23672 17408 23724
rect 17460 23672 17466 23724
rect 17678 23672 17684 23724
rect 17736 23672 17742 23724
rect 24872 23721 24900 23752
rect 25130 23740 25136 23752
rect 25188 23740 25194 23792
rect 26418 23740 26424 23792
rect 26476 23780 26482 23792
rect 38286 23780 38292 23792
rect 26476 23752 38292 23780
rect 26476 23740 26482 23752
rect 38286 23740 38292 23752
rect 38344 23740 38350 23792
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23681 24915 23715
rect 24857 23675 24915 23681
rect 26234 23672 26240 23724
rect 26292 23672 26298 23724
rect 30466 23672 30472 23724
rect 30524 23712 30530 23724
rect 32677 23715 32735 23721
rect 32677 23712 32689 23715
rect 30524 23684 32689 23712
rect 30524 23672 30530 23684
rect 32677 23681 32689 23684
rect 32723 23681 32735 23715
rect 32677 23675 32735 23681
rect 32769 23715 32827 23721
rect 32769 23681 32781 23715
rect 32815 23712 32827 23715
rect 33042 23712 33048 23724
rect 32815 23684 33048 23712
rect 32815 23681 32827 23684
rect 32769 23675 32827 23681
rect 33042 23672 33048 23684
rect 33100 23672 33106 23724
rect 34698 23672 34704 23724
rect 34756 23712 34762 23724
rect 34885 23715 34943 23721
rect 34885 23712 34897 23715
rect 34756 23684 34897 23712
rect 34756 23672 34762 23684
rect 34885 23681 34897 23684
rect 34931 23681 34943 23715
rect 34885 23675 34943 23681
rect 34974 23672 34980 23724
rect 35032 23672 35038 23724
rect 35066 23672 35072 23724
rect 35124 23712 35130 23724
rect 35345 23715 35403 23721
rect 35345 23712 35357 23715
rect 35124 23684 35357 23712
rect 35124 23672 35130 23684
rect 35345 23681 35357 23684
rect 35391 23681 35403 23715
rect 35345 23675 35403 23681
rect 8297 23647 8355 23653
rect 8297 23644 8309 23647
rect 8260 23616 8309 23644
rect 8260 23604 8266 23616
rect 8297 23613 8309 23616
rect 8343 23613 8355 23647
rect 8297 23607 8355 23613
rect 8389 23647 8447 23653
rect 8389 23613 8401 23647
rect 8435 23644 8447 23647
rect 9401 23647 9459 23653
rect 9401 23644 9413 23647
rect 8435 23616 9413 23644
rect 8435 23613 8447 23616
rect 8389 23607 8447 23613
rect 9401 23613 9413 23616
rect 9447 23644 9459 23647
rect 11514 23644 11520 23656
rect 9447 23616 11520 23644
rect 9447 23613 9459 23616
rect 9401 23607 9459 23613
rect 11514 23604 11520 23616
rect 11572 23604 11578 23656
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 14185 23647 14243 23653
rect 14185 23644 14197 23647
rect 12032 23616 14197 23644
rect 12032 23604 12038 23616
rect 14185 23613 14197 23616
rect 14231 23644 14243 23647
rect 15013 23647 15071 23653
rect 15013 23644 15025 23647
rect 14231 23616 15025 23644
rect 14231 23613 14243 23616
rect 14185 23607 14243 23613
rect 15013 23613 15025 23616
rect 15059 23613 15071 23647
rect 15013 23607 15071 23613
rect 24486 23604 24492 23656
rect 24544 23644 24550 23656
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 24544 23616 25145 23644
rect 24544 23604 24550 23616
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 29270 23604 29276 23656
rect 29328 23644 29334 23656
rect 32861 23647 32919 23653
rect 32861 23644 32873 23647
rect 29328 23616 32873 23644
rect 29328 23604 29334 23616
rect 32861 23613 32873 23616
rect 32907 23644 32919 23647
rect 32950 23644 32956 23656
rect 32907 23616 32956 23644
rect 32907 23613 32919 23616
rect 32861 23607 32919 23613
rect 32950 23604 32956 23616
rect 33008 23604 33014 23656
rect 13538 23576 13544 23588
rect 8036 23548 13544 23576
rect 2280 23536 2286 23548
rect 13538 23536 13544 23548
rect 13596 23536 13602 23588
rect 30374 23536 30380 23588
rect 30432 23576 30438 23588
rect 35084 23576 35112 23672
rect 35894 23576 35900 23588
rect 30432 23548 35112 23576
rect 35360 23548 35900 23576
rect 30432 23536 30438 23548
rect 2958 23468 2964 23520
rect 3016 23508 3022 23520
rect 6549 23511 6607 23517
rect 6549 23508 6561 23511
rect 3016 23480 6561 23508
rect 3016 23468 3022 23480
rect 6549 23477 6561 23480
rect 6595 23477 6607 23511
rect 6549 23471 6607 23477
rect 6822 23468 6828 23520
rect 6880 23508 6886 23520
rect 7837 23511 7895 23517
rect 7837 23508 7849 23511
rect 6880 23480 7849 23508
rect 6880 23468 6886 23480
rect 7837 23477 7849 23480
rect 7883 23477 7895 23511
rect 7837 23471 7895 23477
rect 12158 23468 12164 23520
rect 12216 23508 12222 23520
rect 13081 23511 13139 23517
rect 13081 23508 13093 23511
rect 12216 23480 13093 23508
rect 12216 23468 12222 23480
rect 13081 23477 13093 23480
rect 13127 23477 13139 23511
rect 13081 23471 13139 23477
rect 17862 23468 17868 23520
rect 17920 23508 17926 23520
rect 18233 23511 18291 23517
rect 18233 23508 18245 23511
rect 17920 23480 18245 23508
rect 17920 23468 17926 23480
rect 18233 23477 18245 23480
rect 18279 23477 18291 23511
rect 18233 23471 18291 23477
rect 26510 23468 26516 23520
rect 26568 23508 26574 23520
rect 26605 23511 26663 23517
rect 26605 23508 26617 23511
rect 26568 23480 26617 23508
rect 26568 23468 26574 23480
rect 26605 23477 26617 23480
rect 26651 23477 26663 23511
rect 26605 23471 26663 23477
rect 31846 23468 31852 23520
rect 31904 23508 31910 23520
rect 35360 23517 35388 23548
rect 35894 23536 35900 23548
rect 35952 23536 35958 23588
rect 32309 23511 32367 23517
rect 32309 23508 32321 23511
rect 31904 23480 32321 23508
rect 31904 23468 31910 23480
rect 32309 23477 32321 23480
rect 32355 23477 32367 23511
rect 32309 23471 32367 23477
rect 35345 23511 35403 23517
rect 35345 23477 35357 23511
rect 35391 23477 35403 23511
rect 35345 23471 35403 23477
rect 35529 23511 35587 23517
rect 35529 23477 35541 23511
rect 35575 23508 35587 23511
rect 35618 23508 35624 23520
rect 35575 23480 35624 23508
rect 35575 23477 35587 23480
rect 35529 23471 35587 23477
rect 35618 23468 35624 23480
rect 35676 23468 35682 23520
rect 1104 23418 39192 23440
rect 1104 23366 5711 23418
rect 5763 23366 5775 23418
rect 5827 23366 5839 23418
rect 5891 23366 5903 23418
rect 5955 23366 5967 23418
rect 6019 23366 15233 23418
rect 15285 23366 15297 23418
rect 15349 23366 15361 23418
rect 15413 23366 15425 23418
rect 15477 23366 15489 23418
rect 15541 23366 24755 23418
rect 24807 23366 24819 23418
rect 24871 23366 24883 23418
rect 24935 23366 24947 23418
rect 24999 23366 25011 23418
rect 25063 23366 34277 23418
rect 34329 23366 34341 23418
rect 34393 23366 34405 23418
rect 34457 23366 34469 23418
rect 34521 23366 34533 23418
rect 34585 23366 39192 23418
rect 1104 23344 39192 23366
rect 8938 23264 8944 23316
rect 8996 23304 9002 23316
rect 9309 23307 9367 23313
rect 9309 23304 9321 23307
rect 8996 23276 9321 23304
rect 8996 23264 9002 23276
rect 9309 23273 9321 23276
rect 9355 23273 9367 23307
rect 9309 23267 9367 23273
rect 9493 23307 9551 23313
rect 9493 23273 9505 23307
rect 9539 23304 9551 23307
rect 12434 23304 12440 23316
rect 9539 23276 12440 23304
rect 9539 23273 9551 23276
rect 9493 23267 9551 23273
rect 12434 23264 12440 23276
rect 12492 23264 12498 23316
rect 25593 23307 25651 23313
rect 25593 23273 25605 23307
rect 25639 23304 25651 23307
rect 26234 23304 26240 23316
rect 25639 23276 26240 23304
rect 25639 23273 25651 23276
rect 25593 23267 25651 23273
rect 26234 23264 26240 23276
rect 26292 23264 26298 23316
rect 29914 23264 29920 23316
rect 29972 23304 29978 23316
rect 31849 23307 31907 23313
rect 31849 23304 31861 23307
rect 29972 23276 31861 23304
rect 29972 23264 29978 23276
rect 31849 23273 31861 23276
rect 31895 23273 31907 23307
rect 31849 23267 31907 23273
rect 2222 23196 2228 23248
rect 2280 23236 2286 23248
rect 19150 23236 19156 23248
rect 2280 23208 19156 23236
rect 2280 23196 2286 23208
rect 19150 23196 19156 23208
rect 19208 23196 19214 23248
rect 3786 23128 3792 23180
rect 3844 23168 3850 23180
rect 6825 23171 6883 23177
rect 6825 23168 6837 23171
rect 3844 23140 6837 23168
rect 3844 23128 3850 23140
rect 6825 23137 6837 23140
rect 6871 23137 6883 23171
rect 6825 23131 6883 23137
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23100 2283 23103
rect 2869 23103 2927 23109
rect 2869 23100 2881 23103
rect 2271 23072 2881 23100
rect 2271 23069 2283 23072
rect 2225 23063 2283 23069
rect 2869 23069 2881 23072
rect 2915 23100 2927 23103
rect 4062 23100 4068 23112
rect 2915 23072 4068 23100
rect 2915 23069 2927 23072
rect 2869 23063 2927 23069
rect 4062 23060 4068 23072
rect 4120 23060 4126 23112
rect 2317 23035 2375 23041
rect 2317 23001 2329 23035
rect 2363 23032 2375 23035
rect 4706 23032 4712 23044
rect 2363 23004 4712 23032
rect 2363 23001 2375 23004
rect 2317 22995 2375 23001
rect 4706 22992 4712 23004
rect 4764 22992 4770 23044
rect 6840 23032 6868 23131
rect 7006 23128 7012 23180
rect 7064 23168 7070 23180
rect 8110 23168 8116 23180
rect 7064 23140 8116 23168
rect 7064 23128 7070 23140
rect 8110 23128 8116 23140
rect 8168 23128 8174 23180
rect 13538 23128 13544 23180
rect 13596 23128 13602 23180
rect 19242 23168 19248 23180
rect 13648 23140 19248 23168
rect 10689 23103 10747 23109
rect 10689 23069 10701 23103
rect 10735 23100 10747 23103
rect 11882 23100 11888 23112
rect 10735 23072 11888 23100
rect 10735 23069 10747 23072
rect 10689 23063 10747 23069
rect 11882 23060 11888 23072
rect 11940 23100 11946 23112
rect 13648 23100 13676 23140
rect 19242 23128 19248 23140
rect 19300 23128 19306 23180
rect 23937 23171 23995 23177
rect 23937 23137 23949 23171
rect 23983 23168 23995 23171
rect 27890 23168 27896 23180
rect 23983 23140 27896 23168
rect 23983 23137 23995 23140
rect 23937 23131 23995 23137
rect 27890 23128 27896 23140
rect 27948 23128 27954 23180
rect 11940 23072 13676 23100
rect 11940 23060 11946 23072
rect 13722 23060 13728 23112
rect 13780 23100 13786 23112
rect 14277 23103 14335 23109
rect 14277 23100 14289 23103
rect 13780 23072 14289 23100
rect 13780 23060 13786 23072
rect 14277 23069 14289 23072
rect 14323 23100 14335 23103
rect 14826 23100 14832 23112
rect 14323 23072 14832 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 16666 23060 16672 23112
rect 16724 23100 16730 23112
rect 23661 23103 23719 23109
rect 23661 23100 23673 23103
rect 16724 23072 23673 23100
rect 16724 23060 16730 23072
rect 23661 23069 23673 23072
rect 23707 23100 23719 23103
rect 25314 23100 25320 23112
rect 23707 23072 25320 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 25314 23060 25320 23072
rect 25372 23060 25378 23112
rect 25498 23060 25504 23112
rect 25556 23060 25562 23112
rect 9125 23035 9183 23041
rect 9125 23032 9137 23035
rect 6840 23004 9137 23032
rect 9125 23001 9137 23004
rect 9171 23001 9183 23035
rect 9125 22995 9183 23001
rect 11238 22992 11244 23044
rect 11296 22992 11302 23044
rect 13538 23032 13544 23044
rect 13004 23004 13544 23032
rect 2961 22967 3019 22973
rect 2961 22933 2973 22967
rect 3007 22964 3019 22967
rect 3510 22964 3516 22976
rect 3007 22936 3516 22964
rect 3007 22933 3019 22936
rect 2961 22927 3019 22933
rect 3510 22924 3516 22936
rect 3568 22924 3574 22976
rect 6270 22924 6276 22976
rect 6328 22964 6334 22976
rect 6365 22967 6423 22973
rect 6365 22964 6377 22967
rect 6328 22936 6377 22964
rect 6328 22924 6334 22936
rect 6365 22933 6377 22936
rect 6411 22933 6423 22967
rect 6365 22927 6423 22933
rect 6730 22924 6736 22976
rect 6788 22924 6794 22976
rect 9306 22924 9312 22976
rect 9364 22973 9370 22976
rect 13004 22973 13032 23004
rect 13538 22992 13544 23004
rect 13596 22992 13602 23044
rect 18598 22992 18604 23044
rect 18656 23032 18662 23044
rect 26878 23032 26884 23044
rect 18656 23004 26884 23032
rect 18656 22992 18662 23004
rect 26878 22992 26884 23004
rect 26936 22992 26942 23044
rect 31665 23035 31723 23041
rect 31665 23001 31677 23035
rect 31711 23032 31723 23035
rect 33042 23032 33048 23044
rect 31711 23004 33048 23032
rect 31711 23001 31723 23004
rect 31665 22995 31723 23001
rect 33042 22992 33048 23004
rect 33100 22992 33106 23044
rect 9364 22967 9383 22973
rect 9371 22933 9383 22967
rect 9364 22927 9383 22933
rect 12989 22967 13047 22973
rect 12989 22933 13001 22967
rect 13035 22933 13047 22967
rect 12989 22927 13047 22933
rect 9364 22924 9370 22927
rect 13262 22924 13268 22976
rect 13320 22964 13326 22976
rect 13357 22967 13415 22973
rect 13357 22964 13369 22967
rect 13320 22936 13369 22964
rect 13320 22924 13326 22936
rect 13357 22933 13369 22936
rect 13403 22933 13415 22967
rect 13357 22927 13415 22933
rect 13446 22924 13452 22976
rect 13504 22924 13510 22976
rect 14366 22924 14372 22976
rect 14424 22924 14430 22976
rect 22646 22924 22652 22976
rect 22704 22964 22710 22976
rect 23293 22967 23351 22973
rect 23293 22964 23305 22967
rect 22704 22936 23305 22964
rect 22704 22924 22710 22936
rect 23293 22933 23305 22936
rect 23339 22933 23351 22967
rect 23293 22927 23351 22933
rect 23753 22967 23811 22973
rect 23753 22933 23765 22967
rect 23799 22964 23811 22967
rect 24118 22964 24124 22976
rect 23799 22936 24124 22964
rect 23799 22933 23811 22936
rect 23753 22927 23811 22933
rect 24118 22924 24124 22936
rect 24176 22924 24182 22976
rect 30006 22924 30012 22976
rect 30064 22964 30070 22976
rect 31865 22967 31923 22973
rect 31865 22964 31877 22967
rect 30064 22936 31877 22964
rect 30064 22924 30070 22936
rect 31865 22933 31877 22936
rect 31911 22933 31923 22967
rect 31865 22927 31923 22933
rect 32033 22967 32091 22973
rect 32033 22933 32045 22967
rect 32079 22964 32091 22967
rect 32122 22964 32128 22976
rect 32079 22936 32128 22964
rect 32079 22933 32091 22936
rect 32033 22927 32091 22933
rect 32122 22924 32128 22936
rect 32180 22924 32186 22976
rect 1104 22874 39352 22896
rect 1104 22822 10472 22874
rect 10524 22822 10536 22874
rect 10588 22822 10600 22874
rect 10652 22822 10664 22874
rect 10716 22822 10728 22874
rect 10780 22822 19994 22874
rect 20046 22822 20058 22874
rect 20110 22822 20122 22874
rect 20174 22822 20186 22874
rect 20238 22822 20250 22874
rect 20302 22822 29516 22874
rect 29568 22822 29580 22874
rect 29632 22822 29644 22874
rect 29696 22822 29708 22874
rect 29760 22822 29772 22874
rect 29824 22822 39038 22874
rect 39090 22822 39102 22874
rect 39154 22822 39166 22874
rect 39218 22822 39230 22874
rect 39282 22822 39294 22874
rect 39346 22822 39352 22874
rect 1104 22800 39352 22822
rect 2222 22720 2228 22772
rect 2280 22720 2286 22772
rect 4735 22763 4793 22769
rect 4735 22729 4747 22763
rect 4781 22760 4793 22763
rect 9306 22760 9312 22772
rect 4781 22732 9312 22760
rect 4781 22729 4793 22732
rect 4735 22723 4793 22729
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 18782 22760 18788 22772
rect 12406 22732 18788 22760
rect 1673 22695 1731 22701
rect 1673 22661 1685 22695
rect 1719 22692 1731 22695
rect 2240 22692 2268 22720
rect 1719 22664 2268 22692
rect 4525 22695 4583 22701
rect 1719 22661 1731 22664
rect 1673 22655 1731 22661
rect 4525 22661 4537 22695
rect 4571 22661 4583 22695
rect 7650 22692 7656 22704
rect 4525 22655 4583 22661
rect 5736 22664 7656 22692
rect 3605 22627 3663 22633
rect 3605 22593 3617 22627
rect 3651 22624 3663 22627
rect 4062 22624 4068 22636
rect 3651 22596 4068 22624
rect 3651 22593 3663 22596
rect 3605 22587 3663 22593
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 4540 22556 4568 22655
rect 5736 22633 5764 22664
rect 7650 22652 7656 22664
rect 7708 22652 7714 22704
rect 10318 22652 10324 22704
rect 10376 22692 10382 22704
rect 10413 22695 10471 22701
rect 10413 22692 10425 22695
rect 10376 22664 10425 22692
rect 10376 22652 10382 22664
rect 10413 22661 10425 22664
rect 10459 22692 10471 22695
rect 12406 22692 12434 22732
rect 18782 22720 18788 22732
rect 18840 22720 18846 22772
rect 19058 22720 19064 22772
rect 19116 22760 19122 22772
rect 21269 22763 21327 22769
rect 19116 22732 21220 22760
rect 19116 22720 19122 22732
rect 10459 22664 12434 22692
rect 14185 22695 14243 22701
rect 10459 22661 10471 22664
rect 10413 22655 10471 22661
rect 14185 22661 14197 22695
rect 14231 22692 14243 22695
rect 14274 22692 14280 22704
rect 14231 22664 14280 22692
rect 14231 22661 14243 22664
rect 14185 22655 14243 22661
rect 14274 22652 14280 22664
rect 14332 22652 14338 22704
rect 15562 22692 15568 22704
rect 15410 22664 15568 22692
rect 15562 22652 15568 22664
rect 15620 22652 15626 22704
rect 17954 22652 17960 22704
rect 18012 22692 18018 22704
rect 21192 22692 21220 22732
rect 21269 22729 21281 22763
rect 21315 22760 21327 22763
rect 24394 22760 24400 22772
rect 21315 22732 24400 22760
rect 21315 22729 21327 22732
rect 21269 22723 21327 22729
rect 24394 22720 24400 22732
rect 24452 22720 24458 22772
rect 31757 22763 31815 22769
rect 31757 22729 31769 22763
rect 31803 22760 31815 22763
rect 32398 22760 32404 22772
rect 31803 22732 32404 22760
rect 31803 22729 31815 22732
rect 31757 22723 31815 22729
rect 32398 22720 32404 22732
rect 32456 22720 32462 22772
rect 28258 22692 28264 22704
rect 18012 22664 20286 22692
rect 21192 22664 24256 22692
rect 18012 22652 18018 22664
rect 5721 22627 5779 22633
rect 5721 22593 5733 22627
rect 5767 22593 5779 22627
rect 5721 22587 5779 22593
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 10229 22627 10287 22633
rect 5859 22596 9168 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 8202 22556 8208 22568
rect 4540 22528 8208 22556
rect 8202 22516 8208 22528
rect 8260 22556 8266 22568
rect 8846 22556 8852 22568
rect 8260 22528 8852 22556
rect 8260 22516 8266 22528
rect 8846 22516 8852 22528
rect 8904 22516 8910 22568
rect 3970 22448 3976 22500
rect 4028 22488 4034 22500
rect 7006 22488 7012 22500
rect 4028 22460 7012 22488
rect 4028 22448 4034 22460
rect 7006 22448 7012 22460
rect 7064 22448 7070 22500
rect 934 22380 940 22432
rect 992 22420 998 22432
rect 1765 22423 1823 22429
rect 1765 22420 1777 22423
rect 992 22392 1777 22420
rect 992 22380 998 22392
rect 1765 22389 1777 22392
rect 1811 22389 1823 22423
rect 1765 22383 1823 22389
rect 3694 22380 3700 22432
rect 3752 22380 3758 22432
rect 4709 22423 4767 22429
rect 4709 22389 4721 22423
rect 4755 22420 4767 22423
rect 4798 22420 4804 22432
rect 4755 22392 4804 22420
rect 4755 22389 4767 22392
rect 4709 22383 4767 22389
rect 4798 22380 4804 22392
rect 4856 22380 4862 22432
rect 4893 22423 4951 22429
rect 4893 22389 4905 22423
rect 4939 22420 4951 22423
rect 5626 22420 5632 22432
rect 4939 22392 5632 22420
rect 4939 22389 4951 22392
rect 4893 22383 4951 22389
rect 5626 22380 5632 22392
rect 5684 22380 5690 22432
rect 5997 22423 6055 22429
rect 5997 22389 6009 22423
rect 6043 22420 6055 22423
rect 6178 22420 6184 22432
rect 6043 22392 6184 22420
rect 6043 22389 6055 22392
rect 5997 22383 6055 22389
rect 6178 22380 6184 22392
rect 6236 22380 6242 22432
rect 9140 22420 9168 22596
rect 10229 22593 10241 22627
rect 10275 22593 10287 22627
rect 10229 22587 10287 22593
rect 10689 22627 10747 22633
rect 10689 22593 10701 22627
rect 10735 22624 10747 22627
rect 11238 22624 11244 22636
rect 10735 22596 11244 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 10244 22556 10272 22587
rect 11238 22584 11244 22596
rect 11296 22584 11302 22636
rect 12526 22584 12532 22636
rect 12584 22624 12590 22636
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12584 22596 12909 22624
rect 12584 22584 12590 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 13906 22584 13912 22636
rect 13964 22584 13970 22636
rect 18414 22584 18420 22636
rect 18472 22584 18478 22636
rect 11330 22556 11336 22568
rect 10244 22528 11336 22556
rect 11330 22516 11336 22528
rect 11388 22516 11394 22568
rect 13078 22516 13084 22568
rect 13136 22516 13142 22568
rect 14642 22516 14648 22568
rect 14700 22556 14706 22568
rect 15933 22559 15991 22565
rect 15933 22556 15945 22559
rect 14700 22528 15945 22556
rect 14700 22516 14706 22528
rect 15933 22525 15945 22528
rect 15979 22556 15991 22559
rect 15979 22528 16574 22556
rect 15979 22525 15991 22528
rect 15933 22519 15991 22525
rect 16546 22488 16574 22528
rect 18690 22516 18696 22568
rect 18748 22516 18754 22568
rect 19521 22559 19579 22565
rect 19521 22525 19533 22559
rect 19567 22556 19579 22559
rect 19797 22559 19855 22565
rect 19567 22528 19656 22556
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 19334 22488 19340 22500
rect 16546 22460 19340 22488
rect 19334 22448 19340 22460
rect 19392 22448 19398 22500
rect 14550 22420 14556 22432
rect 9140 22392 14556 22420
rect 14550 22380 14556 22392
rect 14608 22380 14614 22432
rect 19628 22420 19656 22528
rect 19797 22525 19809 22559
rect 19843 22556 19855 22559
rect 24228 22556 24256 22664
rect 24320 22664 28264 22692
rect 24320 22633 24348 22664
rect 28258 22652 28264 22664
rect 28316 22652 28322 22704
rect 32309 22695 32367 22701
rect 32309 22661 32321 22695
rect 32355 22692 32367 22695
rect 37090 22692 37096 22704
rect 32355 22664 37096 22692
rect 32355 22661 32367 22664
rect 32309 22655 32367 22661
rect 37090 22652 37096 22664
rect 37148 22652 37154 22704
rect 24305 22627 24363 22633
rect 24305 22593 24317 22627
rect 24351 22593 24363 22627
rect 24305 22587 24363 22593
rect 24394 22584 24400 22636
rect 24452 22624 24458 22636
rect 28994 22624 29000 22636
rect 24452 22596 29000 22624
rect 24452 22584 24458 22596
rect 28994 22584 29000 22596
rect 29052 22584 29058 22636
rect 31386 22584 31392 22636
rect 31444 22584 31450 22636
rect 31573 22627 31631 22633
rect 31573 22593 31585 22627
rect 31619 22624 31631 22627
rect 32950 22624 32956 22636
rect 31619 22596 32956 22624
rect 31619 22593 31631 22596
rect 31573 22587 31631 22593
rect 32950 22584 32956 22596
rect 33008 22584 33014 22636
rect 24581 22559 24639 22565
rect 24581 22556 24593 22559
rect 19843 22528 23980 22556
rect 24228 22528 24593 22556
rect 19843 22525 19855 22528
rect 19797 22519 19855 22525
rect 22278 22488 22284 22500
rect 20824 22460 22284 22488
rect 20824 22420 20852 22460
rect 22278 22448 22284 22460
rect 22336 22448 22342 22500
rect 23952 22497 23980 22528
rect 24581 22525 24593 22528
rect 24627 22556 24639 22559
rect 25222 22556 25228 22568
rect 24627 22528 25228 22556
rect 24627 22525 24639 22528
rect 24581 22519 24639 22525
rect 25222 22516 25228 22528
rect 25280 22516 25286 22568
rect 26878 22516 26884 22568
rect 26936 22556 26942 22568
rect 33045 22559 33103 22565
rect 26936 22528 32996 22556
rect 26936 22516 26942 22528
rect 23937 22491 23995 22497
rect 23937 22457 23949 22491
rect 23983 22457 23995 22491
rect 32122 22488 32128 22500
rect 23937 22451 23995 22457
rect 31588 22460 32128 22488
rect 31588 22429 31616 22460
rect 32122 22448 32128 22460
rect 32180 22448 32186 22500
rect 32968 22488 32996 22528
rect 33045 22525 33057 22559
rect 33091 22556 33103 22559
rect 33134 22556 33140 22568
rect 33091 22528 33140 22556
rect 33091 22525 33103 22528
rect 33045 22519 33103 22525
rect 33134 22516 33140 22528
rect 33192 22516 33198 22568
rect 33962 22488 33968 22500
rect 32968 22460 33968 22488
rect 33962 22448 33968 22460
rect 34020 22448 34026 22500
rect 19628 22392 20852 22420
rect 31573 22423 31631 22429
rect 31573 22389 31585 22423
rect 31619 22389 31631 22423
rect 31573 22383 31631 22389
rect 1104 22330 39192 22352
rect 1104 22278 5711 22330
rect 5763 22278 5775 22330
rect 5827 22278 5839 22330
rect 5891 22278 5903 22330
rect 5955 22278 5967 22330
rect 6019 22278 15233 22330
rect 15285 22278 15297 22330
rect 15349 22278 15361 22330
rect 15413 22278 15425 22330
rect 15477 22278 15489 22330
rect 15541 22278 24755 22330
rect 24807 22278 24819 22330
rect 24871 22278 24883 22330
rect 24935 22278 24947 22330
rect 24999 22278 25011 22330
rect 25063 22278 34277 22330
rect 34329 22278 34341 22330
rect 34393 22278 34405 22330
rect 34457 22278 34469 22330
rect 34521 22278 34533 22330
rect 34585 22278 39192 22330
rect 1104 22256 39192 22278
rect 4798 22176 4804 22228
rect 4856 22216 4862 22228
rect 8938 22216 8944 22228
rect 4856 22188 8944 22216
rect 4856 22176 4862 22188
rect 8938 22176 8944 22188
rect 8996 22176 9002 22228
rect 25222 22176 25228 22228
rect 25280 22216 25286 22228
rect 32582 22216 32588 22228
rect 25280 22188 32588 22216
rect 25280 22176 25286 22188
rect 32582 22176 32588 22188
rect 32640 22176 32646 22228
rect 3970 22148 3976 22160
rect 3436 22120 3976 22148
rect 3436 22094 3464 22120
rect 3970 22108 3976 22120
rect 4028 22108 4034 22160
rect 4890 22148 4896 22160
rect 4724 22120 4896 22148
rect 4724 22094 4752 22120
rect 4890 22108 4896 22120
rect 4948 22108 4954 22160
rect 13630 22148 13636 22160
rect 13556 22120 13636 22148
rect 3344 22092 3464 22094
rect 3326 22080 3332 22092
rect 3287 22052 3332 22080
rect 3326 22040 3332 22052
rect 3384 22066 3464 22092
rect 4632 22089 4752 22094
rect 4617 22083 4752 22089
rect 3384 22040 3390 22066
rect 4617 22049 4629 22083
rect 4663 22066 4752 22083
rect 10689 22083 10747 22089
rect 4663 22052 4697 22066
rect 4663 22049 4675 22052
rect 4617 22043 4675 22049
rect 10689 22049 10701 22083
rect 10735 22080 10747 22083
rect 12434 22080 12440 22092
rect 10735 22052 12440 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 12434 22040 12440 22052
rect 12492 22080 12498 22092
rect 13556 22089 13584 22120
rect 13630 22108 13636 22120
rect 13688 22148 13694 22160
rect 18598 22148 18604 22160
rect 13688 22120 18604 22148
rect 13688 22108 13694 22120
rect 18598 22108 18604 22120
rect 18656 22108 18662 22160
rect 30282 22108 30288 22160
rect 30340 22148 30346 22160
rect 33134 22148 33140 22160
rect 30340 22120 33140 22148
rect 30340 22108 30346 22120
rect 13541 22083 13599 22089
rect 12492 22052 13400 22080
rect 12492 22040 12498 22052
rect 13372 22012 13400 22052
rect 13541 22049 13553 22083
rect 13587 22080 13599 22083
rect 14921 22083 14979 22089
rect 13587 22052 13621 22080
rect 13587 22049 13599 22052
rect 13541 22043 13599 22049
rect 14921 22049 14933 22083
rect 14967 22080 14979 22083
rect 15562 22080 15568 22092
rect 14967 22052 15568 22080
rect 14967 22049 14979 22052
rect 14921 22043 14979 22049
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 16577 22083 16635 22089
rect 16577 22049 16589 22083
rect 16623 22080 16635 22083
rect 17954 22080 17960 22092
rect 16623 22052 17960 22080
rect 16623 22049 16635 22052
rect 16577 22043 16635 22049
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 27706 22040 27712 22092
rect 27764 22080 27770 22092
rect 31478 22080 31484 22092
rect 27764 22052 31484 22080
rect 27764 22040 27770 22052
rect 31478 22040 31484 22052
rect 31536 22080 31542 22092
rect 32968 22089 32996 22120
rect 33134 22108 33140 22120
rect 33192 22108 33198 22160
rect 31573 22083 31631 22089
rect 31573 22080 31585 22083
rect 31536 22052 31585 22080
rect 31536 22040 31542 22052
rect 31573 22049 31585 22052
rect 31619 22049 31631 22083
rect 31573 22043 31631 22049
rect 32953 22083 33011 22089
rect 32953 22049 32965 22083
rect 32999 22080 33011 22083
rect 32999 22052 33033 22080
rect 32999 22049 33011 22052
rect 32953 22043 33011 22049
rect 13906 22012 13912 22024
rect 13372 21984 13912 22012
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14826 21972 14832 22024
rect 14884 22012 14890 22024
rect 15841 22015 15899 22021
rect 15841 22012 15853 22015
rect 14884 21984 15853 22012
rect 14884 21972 14890 21984
rect 15841 21981 15853 21984
rect 15887 22012 15899 22015
rect 16485 22015 16543 22021
rect 16485 22012 16497 22015
rect 15887 21984 16497 22012
rect 15887 21981 15899 21984
rect 15841 21975 15899 21981
rect 16485 21981 16497 21984
rect 16531 22012 16543 22015
rect 18601 22015 18659 22021
rect 18601 22012 18613 22015
rect 16531 21984 18613 22012
rect 16531 21981 16543 21984
rect 16485 21975 16543 21981
rect 18601 21981 18613 21984
rect 18647 22012 18659 22015
rect 18690 22012 18696 22024
rect 18647 21984 18696 22012
rect 18647 21981 18659 21984
rect 18601 21975 18659 21981
rect 18690 21972 18696 21984
rect 18748 21972 18754 22024
rect 26694 22012 26700 22024
rect 22066 21984 26700 22012
rect 4246 21944 4252 21956
rect 2700 21916 4252 21944
rect 2700 21885 2728 21916
rect 4246 21904 4252 21916
rect 4304 21904 4310 21956
rect 10965 21947 11023 21953
rect 10965 21913 10977 21947
rect 11011 21944 11023 21947
rect 11011 21916 11376 21944
rect 11011 21913 11023 21916
rect 10965 21907 11023 21913
rect 2685 21879 2743 21885
rect 2685 21845 2697 21879
rect 2731 21845 2743 21879
rect 2685 21839 2743 21845
rect 3050 21836 3056 21888
rect 3108 21836 3114 21888
rect 3145 21879 3203 21885
rect 3145 21845 3157 21879
rect 3191 21876 3203 21879
rect 3602 21876 3608 21888
rect 3191 21848 3608 21876
rect 3191 21845 3203 21848
rect 3145 21839 3203 21845
rect 3602 21836 3608 21848
rect 3660 21836 3666 21888
rect 3878 21836 3884 21888
rect 3936 21876 3942 21888
rect 3973 21879 4031 21885
rect 3973 21876 3985 21879
rect 3936 21848 3985 21876
rect 3936 21836 3942 21848
rect 3973 21845 3985 21848
rect 4019 21845 4031 21879
rect 3973 21839 4031 21845
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4341 21879 4399 21885
rect 4341 21876 4353 21879
rect 4212 21848 4353 21876
rect 4212 21836 4218 21848
rect 4341 21845 4353 21848
rect 4387 21845 4399 21879
rect 4341 21839 4399 21845
rect 4430 21836 4436 21888
rect 4488 21836 4494 21888
rect 11348 21876 11376 21916
rect 11698 21904 11704 21956
rect 11756 21904 11762 21956
rect 13265 21947 13323 21953
rect 12268 21916 12940 21944
rect 12268 21876 12296 21916
rect 11348 21848 12296 21876
rect 12437 21879 12495 21885
rect 12437 21845 12449 21879
rect 12483 21876 12495 21879
rect 12802 21876 12808 21888
rect 12483 21848 12808 21876
rect 12483 21845 12495 21848
rect 12437 21839 12495 21845
rect 12802 21836 12808 21848
rect 12860 21836 12866 21888
rect 12912 21885 12940 21916
rect 13265 21913 13277 21947
rect 13311 21944 13323 21947
rect 13722 21944 13728 21956
rect 13311 21916 13728 21944
rect 13311 21913 13323 21916
rect 13265 21907 13323 21913
rect 13722 21904 13728 21916
rect 13780 21904 13786 21956
rect 15933 21947 15991 21953
rect 15933 21913 15945 21947
rect 15979 21944 15991 21947
rect 18966 21944 18972 21956
rect 15979 21916 18972 21944
rect 15979 21913 15991 21916
rect 15933 21907 15991 21913
rect 18966 21904 18972 21916
rect 19024 21904 19030 21956
rect 19242 21904 19248 21956
rect 19300 21944 19306 21956
rect 22066 21944 22094 21984
rect 26694 21972 26700 21984
rect 26752 21972 26758 22024
rect 28534 21972 28540 22024
rect 28592 22012 28598 22024
rect 28718 22012 28724 22024
rect 28592 21984 28724 22012
rect 28592 21972 28598 21984
rect 28718 21972 28724 21984
rect 28776 21972 28782 22024
rect 30193 22015 30251 22021
rect 30193 21981 30205 22015
rect 30239 22012 30251 22015
rect 31018 22012 31024 22024
rect 30239 21984 31024 22012
rect 30239 21981 30251 21984
rect 30193 21975 30251 21981
rect 31018 21972 31024 21984
rect 31076 21972 31082 22024
rect 31294 21972 31300 22024
rect 31352 21972 31358 22024
rect 31588 21984 31754 22012
rect 19300 21916 22094 21944
rect 19300 21904 19306 21916
rect 25038 21904 25044 21956
rect 25096 21944 25102 21956
rect 31588 21944 31616 21984
rect 25096 21916 31616 21944
rect 31726 21944 31754 21984
rect 31726 21916 32444 21944
rect 25096 21904 25102 21916
rect 12897 21879 12955 21885
rect 12897 21845 12909 21879
rect 12943 21845 12955 21879
rect 12897 21839 12955 21845
rect 12986 21836 12992 21888
rect 13044 21876 13050 21888
rect 13354 21876 13360 21888
rect 13044 21848 13360 21876
rect 13044 21836 13050 21848
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 18690 21836 18696 21888
rect 18748 21836 18754 21888
rect 28626 21836 28632 21888
rect 28684 21836 28690 21888
rect 29086 21836 29092 21888
rect 29144 21876 29150 21888
rect 32416 21885 32444 21916
rect 30285 21879 30343 21885
rect 30285 21876 30297 21879
rect 29144 21848 30297 21876
rect 29144 21836 29150 21848
rect 30285 21845 30297 21848
rect 30331 21845 30343 21879
rect 30285 21839 30343 21845
rect 32401 21879 32459 21885
rect 32401 21845 32413 21879
rect 32447 21845 32459 21879
rect 32401 21839 32459 21845
rect 32766 21836 32772 21888
rect 32824 21836 32830 21888
rect 32858 21836 32864 21888
rect 32916 21836 32922 21888
rect 1104 21786 39352 21808
rect 1104 21734 10472 21786
rect 10524 21734 10536 21786
rect 10588 21734 10600 21786
rect 10652 21734 10664 21786
rect 10716 21734 10728 21786
rect 10780 21734 19994 21786
rect 20046 21734 20058 21786
rect 20110 21734 20122 21786
rect 20174 21734 20186 21786
rect 20238 21734 20250 21786
rect 20302 21734 29516 21786
rect 29568 21734 29580 21786
rect 29632 21734 29644 21786
rect 29696 21734 29708 21786
rect 29760 21734 29772 21786
rect 29824 21734 39038 21786
rect 39090 21734 39102 21786
rect 39154 21734 39166 21786
rect 39218 21734 39230 21786
rect 39282 21734 39294 21786
rect 39346 21734 39352 21786
rect 1104 21712 39352 21734
rect 4062 21632 4068 21684
rect 4120 21632 4126 21684
rect 4430 21632 4436 21684
rect 4488 21672 4494 21684
rect 11974 21672 11980 21684
rect 4488 21644 11980 21672
rect 4488 21632 4494 21644
rect 11974 21632 11980 21644
rect 12032 21632 12038 21684
rect 13173 21675 13231 21681
rect 13173 21641 13185 21675
rect 13219 21672 13231 21675
rect 15838 21672 15844 21684
rect 13219 21644 15844 21672
rect 13219 21641 13231 21644
rect 13173 21635 13231 21641
rect 15838 21632 15844 21644
rect 15896 21632 15902 21684
rect 16758 21632 16764 21684
rect 16816 21672 16822 21684
rect 26513 21675 26571 21681
rect 16816 21644 17356 21672
rect 16816 21632 16822 21644
rect 12897 21607 12955 21613
rect 12897 21573 12909 21607
rect 12943 21573 12955 21607
rect 12897 21567 12955 21573
rect 3973 21539 4031 21545
rect 3973 21505 3985 21539
rect 4019 21536 4031 21539
rect 4522 21536 4528 21548
rect 4019 21508 4528 21536
rect 4019 21505 4031 21508
rect 3973 21499 4031 21505
rect 4522 21496 4528 21508
rect 4580 21496 4586 21548
rect 12618 21496 12624 21548
rect 12676 21496 12682 21548
rect 12802 21496 12808 21548
rect 12860 21496 12866 21548
rect 12912 21468 12940 21567
rect 17218 21564 17224 21616
rect 17276 21564 17282 21616
rect 17328 21604 17356 21644
rect 26513 21641 26525 21675
rect 26559 21672 26571 21675
rect 27614 21672 27620 21684
rect 26559 21644 27620 21672
rect 26559 21641 26571 21644
rect 26513 21635 26571 21641
rect 27614 21632 27620 21644
rect 27672 21632 27678 21684
rect 31754 21672 31760 21684
rect 28276 21644 31760 21672
rect 25130 21604 25136 21616
rect 17328 21576 17710 21604
rect 24780 21576 25136 21604
rect 13013 21539 13071 21545
rect 13013 21505 13025 21539
rect 13059 21536 13071 21539
rect 13170 21536 13176 21548
rect 13059 21508 13176 21536
rect 13059 21505 13071 21508
rect 13013 21499 13071 21505
rect 13170 21496 13176 21508
rect 13228 21536 13234 21548
rect 24780 21545 24808 21576
rect 25130 21564 25136 21576
rect 25188 21564 25194 21616
rect 28276 21545 28304 21644
rect 31754 21632 31760 21644
rect 31812 21632 31818 21684
rect 28626 21564 28632 21616
rect 28684 21604 28690 21616
rect 31205 21607 31263 21613
rect 28684 21576 29026 21604
rect 28684 21564 28690 21576
rect 31205 21573 31217 21607
rect 31251 21604 31263 21607
rect 31386 21604 31392 21616
rect 31251 21576 31392 21604
rect 31251 21573 31263 21576
rect 31205 21567 31263 21573
rect 31386 21564 31392 21576
rect 31444 21564 31450 21616
rect 24765 21539 24823 21545
rect 13228 21508 15148 21536
rect 13228 21496 13234 21508
rect 13262 21468 13268 21480
rect 12912 21440 13268 21468
rect 13262 21428 13268 21440
rect 13320 21468 13326 21480
rect 15010 21468 15016 21480
rect 13320 21440 15016 21468
rect 13320 21428 13326 21440
rect 15010 21428 15016 21440
rect 15068 21428 15074 21480
rect 15120 21400 15148 21508
rect 24765 21505 24777 21539
rect 24811 21505 24823 21539
rect 28261 21539 28319 21545
rect 24765 21499 24823 21505
rect 16850 21428 16856 21480
rect 16908 21468 16914 21480
rect 16945 21471 17003 21477
rect 16945 21468 16957 21471
rect 16908 21440 16957 21468
rect 16908 21428 16914 21440
rect 16945 21437 16957 21440
rect 16991 21437 17003 21471
rect 16945 21431 17003 21437
rect 17052 21440 18276 21468
rect 17052 21400 17080 21440
rect 15120 21372 17080 21400
rect 18248 21400 18276 21440
rect 18966 21428 18972 21480
rect 19024 21468 19030 21480
rect 23474 21468 23480 21480
rect 19024 21440 23480 21468
rect 19024 21428 19030 21440
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 25038 21428 25044 21480
rect 25096 21428 25102 21480
rect 19702 21400 19708 21412
rect 18248 21372 19708 21400
rect 19702 21360 19708 21372
rect 19760 21360 19766 21412
rect 26160 21400 26188 21522
rect 28261 21505 28273 21539
rect 28307 21505 28319 21539
rect 28261 21499 28319 21505
rect 31018 21496 31024 21548
rect 31076 21536 31082 21548
rect 35713 21539 35771 21545
rect 35713 21536 35725 21539
rect 31076 21508 35725 21536
rect 31076 21496 31082 21508
rect 35713 21505 35725 21508
rect 35759 21536 35771 21539
rect 36078 21536 36084 21548
rect 35759 21508 36084 21536
rect 35759 21505 35771 21508
rect 35713 21499 35771 21505
rect 36078 21496 36084 21508
rect 36136 21536 36142 21548
rect 37550 21536 37556 21548
rect 36136 21508 37556 21536
rect 36136 21496 36142 21508
rect 37550 21496 37556 21508
rect 37608 21496 37614 21548
rect 28534 21428 28540 21480
rect 28592 21428 28598 21480
rect 31294 21428 31300 21480
rect 31352 21428 31358 21480
rect 31478 21428 31484 21480
rect 31536 21428 31542 21480
rect 35805 21403 35863 21409
rect 35805 21400 35817 21403
rect 26160 21372 28396 21400
rect 12618 21292 12624 21344
rect 12676 21332 12682 21344
rect 18693 21335 18751 21341
rect 18693 21332 18705 21335
rect 12676 21304 18705 21332
rect 12676 21292 12682 21304
rect 18693 21301 18705 21304
rect 18739 21301 18751 21335
rect 28368 21332 28396 21372
rect 29564 21372 35817 21400
rect 29564 21332 29592 21372
rect 35805 21369 35817 21372
rect 35851 21369 35863 21403
rect 35805 21363 35863 21369
rect 28368 21304 29592 21332
rect 18693 21295 18751 21301
rect 30006 21292 30012 21344
rect 30064 21292 30070 21344
rect 30834 21292 30840 21344
rect 30892 21292 30898 21344
rect 1104 21242 39192 21264
rect 1104 21190 5711 21242
rect 5763 21190 5775 21242
rect 5827 21190 5839 21242
rect 5891 21190 5903 21242
rect 5955 21190 5967 21242
rect 6019 21190 15233 21242
rect 15285 21190 15297 21242
rect 15349 21190 15361 21242
rect 15413 21190 15425 21242
rect 15477 21190 15489 21242
rect 15541 21190 24755 21242
rect 24807 21190 24819 21242
rect 24871 21190 24883 21242
rect 24935 21190 24947 21242
rect 24999 21190 25011 21242
rect 25063 21190 34277 21242
rect 34329 21190 34341 21242
rect 34393 21190 34405 21242
rect 34457 21190 34469 21242
rect 34521 21190 34533 21242
rect 34585 21190 39192 21242
rect 1104 21168 39192 21190
rect 12526 21088 12532 21140
rect 12584 21128 12590 21140
rect 12802 21128 12808 21140
rect 12584 21100 12808 21128
rect 12584 21088 12590 21100
rect 12802 21088 12808 21100
rect 12860 21088 12866 21140
rect 23658 21088 23664 21140
rect 23716 21128 23722 21140
rect 23716 21100 26464 21128
rect 23716 21088 23722 21100
rect 3050 21020 3056 21072
rect 3108 21060 3114 21072
rect 13722 21060 13728 21072
rect 3108 21032 13728 21060
rect 3108 21020 3114 21032
rect 13722 21020 13728 21032
rect 13780 21060 13786 21072
rect 23566 21060 23572 21072
rect 13780 21032 23572 21060
rect 13780 21020 13786 21032
rect 23566 21020 23572 21032
rect 23624 21020 23630 21072
rect 26436 21060 26464 21100
rect 27798 21088 27804 21140
rect 27856 21088 27862 21140
rect 28718 21128 28724 21140
rect 27908 21100 28724 21128
rect 27908 21060 27936 21100
rect 28718 21088 28724 21100
rect 28776 21088 28782 21140
rect 29822 21088 29828 21140
rect 29880 21128 29886 21140
rect 29917 21131 29975 21137
rect 29917 21128 29929 21131
rect 29880 21100 29929 21128
rect 29880 21088 29886 21100
rect 29917 21097 29929 21100
rect 29963 21128 29975 21131
rect 30190 21128 30196 21140
rect 29963 21100 30196 21128
rect 29963 21097 29975 21100
rect 29917 21091 29975 21097
rect 30190 21088 30196 21100
rect 30248 21088 30254 21140
rect 30834 21060 30840 21072
rect 26436 21032 27936 21060
rect 28092 21032 30840 21060
rect 6362 20952 6368 21004
rect 6420 20992 6426 21004
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 6420 20964 11161 20992
rect 6420 20952 6426 20964
rect 11149 20961 11161 20964
rect 11195 20992 11207 20995
rect 12618 20992 12624 21004
rect 11195 20964 12624 20992
rect 11195 20961 11207 20964
rect 11149 20955 11207 20961
rect 12618 20952 12624 20964
rect 12676 20992 12682 21004
rect 13630 20992 13636 21004
rect 12676 20964 13636 20992
rect 12676 20952 12682 20964
rect 13630 20952 13636 20964
rect 13688 20952 13694 21004
rect 24578 20952 24584 21004
rect 24636 20992 24642 21004
rect 25130 20992 25136 21004
rect 24636 20964 25136 20992
rect 24636 20952 24642 20964
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 25409 20995 25467 21001
rect 25409 20961 25421 20995
rect 25455 20992 25467 20995
rect 28092 20992 28120 21032
rect 30834 21020 30840 21032
rect 30892 21020 30898 21072
rect 25455 20964 28120 20992
rect 25455 20961 25467 20964
rect 25409 20955 25467 20961
rect 28166 20952 28172 21004
rect 28224 20992 28230 21004
rect 28353 20995 28411 21001
rect 28353 20992 28365 20995
rect 28224 20964 28365 20992
rect 28224 20952 28230 20964
rect 28353 20961 28365 20964
rect 28399 20961 28411 20995
rect 31386 20992 31392 21004
rect 28353 20955 28411 20961
rect 29840 20964 31392 20992
rect 934 20884 940 20936
rect 992 20924 998 20936
rect 1581 20927 1639 20933
rect 1581 20924 1593 20927
rect 992 20896 1593 20924
rect 992 20884 998 20896
rect 1581 20893 1593 20896
rect 1627 20893 1639 20927
rect 1581 20887 1639 20893
rect 3973 20927 4031 20933
rect 3973 20893 3985 20927
rect 4019 20924 4031 20927
rect 4062 20924 4068 20936
rect 4019 20896 4068 20924
rect 4019 20893 4031 20896
rect 3973 20887 4031 20893
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20924 12495 20927
rect 12526 20924 12532 20936
rect 12483 20896 12532 20924
rect 12483 20893 12495 20896
rect 12437 20887 12495 20893
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 13262 20884 13268 20936
rect 13320 20884 13326 20936
rect 13725 20927 13783 20933
rect 13725 20893 13737 20927
rect 13771 20924 13783 20927
rect 16666 20924 16672 20936
rect 13771 20896 16672 20924
rect 13771 20893 13783 20896
rect 13725 20887 13783 20893
rect 1857 20859 1915 20865
rect 1857 20825 1869 20859
rect 1903 20856 1915 20859
rect 5534 20856 5540 20868
rect 1903 20828 5540 20856
rect 1903 20825 1915 20828
rect 1857 20819 1915 20825
rect 5534 20816 5540 20828
rect 5592 20816 5598 20868
rect 10318 20816 10324 20868
rect 10376 20856 10382 20868
rect 11057 20859 11115 20865
rect 11057 20856 11069 20859
rect 10376 20828 11069 20856
rect 10376 20816 10382 20828
rect 11057 20825 11069 20828
rect 11103 20825 11115 20859
rect 11057 20819 11115 20825
rect 12894 20816 12900 20868
rect 12952 20816 12958 20868
rect 12986 20816 12992 20868
rect 13044 20856 13050 20868
rect 13740 20856 13768 20887
rect 16666 20884 16672 20896
rect 16724 20884 16730 20936
rect 27798 20924 27804 20936
rect 26542 20896 27804 20924
rect 27798 20884 27804 20896
rect 27856 20884 27862 20936
rect 29840 20924 29868 20964
rect 31386 20952 31392 20964
rect 31444 20952 31450 21004
rect 33686 20952 33692 21004
rect 33744 20992 33750 21004
rect 36909 20995 36967 21001
rect 36909 20992 36921 20995
rect 33744 20964 36921 20992
rect 33744 20952 33750 20964
rect 36909 20961 36921 20964
rect 36955 20961 36967 20995
rect 36909 20955 36967 20961
rect 28092 20896 29868 20924
rect 13044 20828 13768 20856
rect 13044 20816 13050 20828
rect 3970 20748 3976 20800
rect 4028 20788 4034 20800
rect 4065 20791 4123 20797
rect 4065 20788 4077 20791
rect 4028 20760 4077 20788
rect 4028 20748 4034 20760
rect 4065 20757 4077 20760
rect 4111 20757 4123 20791
rect 4065 20751 4123 20757
rect 9858 20748 9864 20800
rect 9916 20788 9922 20800
rect 10597 20791 10655 20797
rect 10597 20788 10609 20791
rect 9916 20760 10609 20788
rect 9916 20748 9922 20760
rect 10597 20757 10609 20760
rect 10643 20757 10655 20791
rect 10597 20751 10655 20757
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 13446 20788 13452 20800
rect 11020 20760 13452 20788
rect 11020 20748 11026 20760
rect 13446 20748 13452 20760
rect 13504 20748 13510 20800
rect 23566 20748 23572 20800
rect 23624 20788 23630 20800
rect 25590 20788 25596 20800
rect 23624 20760 25596 20788
rect 23624 20748 23630 20760
rect 25590 20748 25596 20760
rect 25648 20748 25654 20800
rect 26881 20791 26939 20797
rect 26881 20757 26893 20791
rect 26927 20788 26939 20791
rect 28092 20788 28120 20896
rect 30098 20884 30104 20936
rect 30156 20924 30162 20936
rect 31018 20924 31024 20936
rect 30156 20896 31024 20924
rect 30156 20884 30162 20896
rect 31018 20884 31024 20896
rect 31076 20884 31082 20936
rect 31754 20884 31760 20936
rect 31812 20924 31818 20936
rect 34885 20927 34943 20933
rect 34885 20924 34897 20927
rect 31812 20896 34897 20924
rect 31812 20884 31818 20896
rect 34885 20893 34897 20896
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 28442 20856 28448 20868
rect 28184 20828 28448 20856
rect 28184 20800 28212 20828
rect 28442 20816 28448 20828
rect 28500 20816 28506 20868
rect 28994 20816 29000 20868
rect 29052 20856 29058 20868
rect 29733 20859 29791 20865
rect 29733 20856 29745 20859
rect 29052 20828 29745 20856
rect 29052 20816 29058 20828
rect 29733 20825 29745 20828
rect 29779 20825 29791 20859
rect 32858 20856 32864 20868
rect 29733 20819 29791 20825
rect 30116 20828 32864 20856
rect 26927 20760 28120 20788
rect 26927 20757 26939 20760
rect 26881 20751 26939 20757
rect 28166 20748 28172 20800
rect 28224 20748 28230 20800
rect 28258 20748 28264 20800
rect 28316 20788 28322 20800
rect 28902 20788 28908 20800
rect 28316 20760 28908 20788
rect 28316 20748 28322 20760
rect 28902 20748 28908 20760
rect 28960 20748 28966 20800
rect 29362 20748 29368 20800
rect 29420 20788 29426 20800
rect 29914 20788 29920 20800
rect 29972 20797 29978 20800
rect 30116 20797 30144 20828
rect 32858 20816 32864 20828
rect 32916 20816 32922 20868
rect 35158 20816 35164 20868
rect 35216 20816 35222 20868
rect 36170 20816 36176 20868
rect 36228 20816 36234 20868
rect 38470 20816 38476 20868
rect 38528 20816 38534 20868
rect 38657 20859 38715 20865
rect 38657 20825 38669 20859
rect 38703 20856 38715 20859
rect 39390 20856 39396 20868
rect 38703 20828 39396 20856
rect 38703 20825 38715 20828
rect 38657 20819 38715 20825
rect 39390 20816 39396 20828
rect 39448 20816 39454 20868
rect 29972 20791 29991 20797
rect 29420 20760 29920 20788
rect 29420 20748 29426 20760
rect 29914 20748 29920 20760
rect 29979 20757 29991 20791
rect 29972 20751 29991 20757
rect 30101 20791 30159 20797
rect 30101 20757 30113 20791
rect 30147 20757 30159 20791
rect 30101 20751 30159 20757
rect 29972 20748 29978 20751
rect 30926 20748 30932 20800
rect 30984 20788 30990 20800
rect 31113 20791 31171 20797
rect 31113 20788 31125 20791
rect 30984 20760 31125 20788
rect 30984 20748 30990 20760
rect 31113 20757 31125 20760
rect 31159 20757 31171 20791
rect 31113 20751 31171 20757
rect 1104 20698 39352 20720
rect 1104 20646 10472 20698
rect 10524 20646 10536 20698
rect 10588 20646 10600 20698
rect 10652 20646 10664 20698
rect 10716 20646 10728 20698
rect 10780 20646 19994 20698
rect 20046 20646 20058 20698
rect 20110 20646 20122 20698
rect 20174 20646 20186 20698
rect 20238 20646 20250 20698
rect 20302 20646 29516 20698
rect 29568 20646 29580 20698
rect 29632 20646 29644 20698
rect 29696 20646 29708 20698
rect 29760 20646 29772 20698
rect 29824 20646 39038 20698
rect 39090 20646 39102 20698
rect 39154 20646 39166 20698
rect 39218 20646 39230 20698
rect 39282 20646 39294 20698
rect 39346 20646 39352 20698
rect 1104 20624 39352 20646
rect 11974 20544 11980 20596
rect 12032 20584 12038 20596
rect 14918 20584 14924 20596
rect 12032 20556 14924 20584
rect 12032 20544 12038 20556
rect 14918 20544 14924 20556
rect 14976 20584 14982 20596
rect 15562 20584 15568 20596
rect 14976 20556 15568 20584
rect 14976 20544 14982 20556
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 19794 20544 19800 20596
rect 19852 20584 19858 20596
rect 25406 20584 25412 20596
rect 19852 20556 25412 20584
rect 19852 20544 19858 20556
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 26878 20544 26884 20596
rect 26936 20584 26942 20596
rect 27525 20587 27583 20593
rect 27525 20584 27537 20587
rect 26936 20556 27537 20584
rect 26936 20544 26942 20556
rect 27525 20553 27537 20556
rect 27571 20553 27583 20587
rect 27525 20547 27583 20553
rect 28534 20544 28540 20596
rect 28592 20584 28598 20596
rect 28721 20587 28779 20593
rect 28721 20584 28733 20587
rect 28592 20556 28733 20584
rect 28592 20544 28598 20556
rect 28721 20553 28733 20556
rect 28767 20553 28779 20587
rect 28721 20547 28779 20553
rect 33137 20587 33195 20593
rect 33137 20553 33149 20587
rect 33183 20584 33195 20587
rect 35158 20584 35164 20596
rect 33183 20556 35164 20584
rect 33183 20553 33195 20556
rect 33137 20547 33195 20553
rect 35158 20544 35164 20556
rect 35216 20544 35222 20596
rect 36170 20544 36176 20596
rect 36228 20544 36234 20596
rect 4617 20519 4675 20525
rect 4617 20516 4629 20519
rect 3726 20488 4629 20516
rect 4617 20485 4629 20488
rect 4663 20485 4675 20519
rect 4617 20479 4675 20485
rect 12115 20519 12173 20525
rect 12115 20485 12127 20519
rect 12161 20516 12173 20519
rect 12526 20516 12532 20528
rect 12161 20488 12532 20516
rect 12161 20485 12173 20488
rect 12115 20479 12173 20485
rect 12526 20476 12532 20488
rect 12584 20476 12590 20528
rect 12618 20476 12624 20528
rect 12676 20516 12682 20528
rect 12894 20516 12900 20528
rect 12676 20488 12900 20516
rect 12676 20476 12682 20488
rect 12894 20476 12900 20488
rect 12952 20516 12958 20528
rect 12952 20488 21956 20516
rect 12952 20476 12958 20488
rect 4525 20451 4583 20457
rect 4525 20417 4537 20451
rect 4571 20448 4583 20451
rect 6546 20448 6552 20460
rect 4571 20420 6552 20448
rect 4571 20417 4583 20420
rect 4525 20411 4583 20417
rect 6546 20408 6552 20420
rect 6604 20408 6610 20460
rect 11330 20408 11336 20460
rect 11388 20448 11394 20460
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 11388 20420 11713 20448
rect 11388 20408 11394 20420
rect 11701 20417 11713 20420
rect 11747 20448 11759 20451
rect 12544 20448 12572 20476
rect 21928 20460 21956 20488
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 29181 20519 29239 20525
rect 29181 20516 29193 20519
rect 22152 20488 29193 20516
rect 22152 20476 22158 20488
rect 29181 20485 29193 20488
rect 29227 20516 29239 20519
rect 30006 20516 30012 20528
rect 29227 20488 30012 20516
rect 29227 20485 29239 20488
rect 29181 20479 29239 20485
rect 30006 20476 30012 20488
rect 30064 20476 30070 20528
rect 33597 20519 33655 20525
rect 33597 20485 33609 20519
rect 33643 20516 33655 20519
rect 33686 20516 33692 20528
rect 33643 20488 33692 20516
rect 33643 20485 33655 20488
rect 33597 20479 33655 20485
rect 33686 20476 33692 20488
rect 33744 20476 33750 20528
rect 16942 20448 16948 20460
rect 11747 20420 12020 20448
rect 12544 20420 16948 20448
rect 11747 20417 11759 20420
rect 11701 20411 11759 20417
rect 11992 20392 12020 20420
rect 16942 20408 16948 20420
rect 17000 20448 17006 20460
rect 21177 20451 21235 20457
rect 17000 20420 17448 20448
rect 17000 20408 17006 20420
rect 17420 20392 17448 20420
rect 21177 20417 21189 20451
rect 21223 20448 21235 20451
rect 21266 20448 21272 20460
rect 21223 20420 21272 20448
rect 21223 20417 21235 20420
rect 21177 20411 21235 20417
rect 21266 20408 21272 20420
rect 21324 20408 21330 20460
rect 21910 20408 21916 20460
rect 21968 20448 21974 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21968 20420 22017 20448
rect 21968 20408 21974 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22741 20451 22799 20457
rect 22741 20417 22753 20451
rect 22787 20417 22799 20451
rect 22741 20411 22799 20417
rect 2222 20340 2228 20392
rect 2280 20340 2286 20392
rect 2501 20383 2559 20389
rect 2501 20349 2513 20383
rect 2547 20380 2559 20383
rect 3878 20380 3884 20392
rect 2547 20352 3884 20380
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 3878 20340 3884 20352
rect 3936 20340 3942 20392
rect 11974 20340 11980 20392
rect 12032 20380 12038 20392
rect 13262 20380 13268 20392
rect 12032 20352 13268 20380
rect 12032 20340 12038 20352
rect 13262 20340 13268 20352
rect 13320 20340 13326 20392
rect 17402 20340 17408 20392
rect 17460 20380 17466 20392
rect 21726 20380 21732 20392
rect 17460 20352 21732 20380
rect 17460 20340 17466 20352
rect 21726 20340 21732 20352
rect 21784 20340 21790 20392
rect 22756 20380 22784 20411
rect 23658 20408 23664 20460
rect 23716 20408 23722 20460
rect 23842 20408 23848 20460
rect 23900 20448 23906 20460
rect 29089 20451 29147 20457
rect 29089 20448 29101 20451
rect 23900 20420 29101 20448
rect 23900 20408 23906 20420
rect 29089 20417 29101 20420
rect 29135 20417 29147 20451
rect 29089 20411 29147 20417
rect 32582 20408 32588 20460
rect 32640 20448 32646 20460
rect 33505 20451 33563 20457
rect 33505 20448 33517 20451
rect 32640 20420 33517 20448
rect 32640 20408 32646 20420
rect 33505 20417 33517 20420
rect 33551 20417 33563 20451
rect 33505 20411 33563 20417
rect 36078 20408 36084 20460
rect 36136 20408 36142 20460
rect 23290 20380 23296 20392
rect 22756 20352 23296 20380
rect 23290 20340 23296 20352
rect 23348 20380 23354 20392
rect 25498 20380 25504 20392
rect 23348 20352 25504 20380
rect 23348 20340 23354 20352
rect 25498 20340 25504 20352
rect 25556 20340 25562 20392
rect 27522 20340 27528 20392
rect 27580 20380 27586 20392
rect 27617 20383 27675 20389
rect 27617 20380 27629 20383
rect 27580 20352 27629 20380
rect 27580 20340 27586 20352
rect 27617 20349 27629 20352
rect 27663 20349 27675 20383
rect 27617 20343 27675 20349
rect 27709 20383 27767 20389
rect 27709 20349 27721 20383
rect 27755 20349 27767 20383
rect 27709 20343 27767 20349
rect 29365 20383 29423 20389
rect 29365 20349 29377 20383
rect 29411 20380 29423 20383
rect 29914 20380 29920 20392
rect 29411 20352 29920 20380
rect 29411 20349 29423 20352
rect 29365 20343 29423 20349
rect 12253 20315 12311 20321
rect 12253 20281 12265 20315
rect 12299 20312 12311 20315
rect 12802 20312 12808 20324
rect 12299 20284 12808 20312
rect 12299 20281 12311 20284
rect 12253 20275 12311 20281
rect 12802 20272 12808 20284
rect 12860 20312 12866 20324
rect 13722 20312 13728 20324
rect 12860 20284 13728 20312
rect 12860 20272 12866 20284
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 21082 20272 21088 20324
rect 21140 20312 21146 20324
rect 22189 20315 22247 20321
rect 22189 20312 22201 20315
rect 21140 20284 22201 20312
rect 21140 20272 21146 20284
rect 22189 20281 22201 20284
rect 22235 20312 22247 20315
rect 22235 20284 25084 20312
rect 22235 20281 22247 20284
rect 22189 20275 22247 20281
rect 3973 20247 4031 20253
rect 3973 20213 3985 20247
rect 4019 20244 4031 20247
rect 4154 20244 4160 20256
rect 4019 20216 4160 20244
rect 4019 20213 4031 20216
rect 3973 20207 4031 20213
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 12069 20247 12127 20253
rect 12069 20213 12081 20247
rect 12115 20244 12127 20247
rect 12986 20244 12992 20256
rect 12115 20216 12992 20244
rect 12115 20213 12127 20216
rect 12069 20207 12127 20213
rect 12986 20204 12992 20216
rect 13044 20204 13050 20256
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 14918 20244 14924 20256
rect 13136 20216 14924 20244
rect 13136 20204 13142 20216
rect 14918 20204 14924 20216
rect 14976 20204 14982 20256
rect 18782 20204 18788 20256
rect 18840 20244 18846 20256
rect 21174 20244 21180 20256
rect 18840 20216 21180 20244
rect 18840 20204 18846 20216
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 21361 20247 21419 20253
rect 21361 20213 21373 20247
rect 21407 20244 21419 20247
rect 22370 20244 22376 20256
rect 21407 20216 22376 20244
rect 21407 20213 21419 20216
rect 21361 20207 21419 20213
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 22833 20247 22891 20253
rect 22833 20213 22845 20247
rect 22879 20244 22891 20247
rect 23106 20244 23112 20256
rect 22879 20216 23112 20244
rect 22879 20213 22891 20216
rect 22833 20207 22891 20213
rect 23106 20204 23112 20216
rect 23164 20204 23170 20256
rect 23658 20204 23664 20256
rect 23716 20244 23722 20256
rect 23753 20247 23811 20253
rect 23753 20244 23765 20247
rect 23716 20216 23765 20244
rect 23716 20204 23722 20216
rect 23753 20213 23765 20216
rect 23799 20213 23811 20247
rect 25056 20244 25084 20284
rect 25130 20272 25136 20324
rect 25188 20312 25194 20324
rect 27724 20312 27752 20343
rect 29914 20340 29920 20352
rect 29972 20380 29978 20392
rect 30282 20380 30288 20392
rect 29972 20352 30288 20380
rect 29972 20340 29978 20352
rect 30282 20340 30288 20352
rect 30340 20340 30346 20392
rect 32674 20340 32680 20392
rect 32732 20380 32738 20392
rect 33781 20383 33839 20389
rect 33781 20380 33793 20383
rect 32732 20352 33793 20380
rect 32732 20340 32738 20352
rect 33781 20349 33793 20352
rect 33827 20380 33839 20383
rect 34790 20380 34796 20392
rect 33827 20352 34796 20380
rect 33827 20349 33839 20352
rect 33781 20343 33839 20349
rect 34790 20340 34796 20352
rect 34848 20340 34854 20392
rect 25188 20284 27752 20312
rect 25188 20272 25194 20284
rect 25958 20244 25964 20256
rect 25056 20216 25964 20244
rect 23753 20207 23811 20213
rect 25958 20204 25964 20216
rect 26016 20204 26022 20256
rect 27154 20204 27160 20256
rect 27212 20204 27218 20256
rect 1104 20154 39192 20176
rect 1104 20102 5711 20154
rect 5763 20102 5775 20154
rect 5827 20102 5839 20154
rect 5891 20102 5903 20154
rect 5955 20102 5967 20154
rect 6019 20102 15233 20154
rect 15285 20102 15297 20154
rect 15349 20102 15361 20154
rect 15413 20102 15425 20154
rect 15477 20102 15489 20154
rect 15541 20102 24755 20154
rect 24807 20102 24819 20154
rect 24871 20102 24883 20154
rect 24935 20102 24947 20154
rect 24999 20102 25011 20154
rect 25063 20102 34277 20154
rect 34329 20102 34341 20154
rect 34393 20102 34405 20154
rect 34457 20102 34469 20154
rect 34521 20102 34533 20154
rect 34585 20102 39192 20154
rect 1104 20080 39192 20102
rect 5994 20000 6000 20052
rect 6052 20000 6058 20052
rect 11330 20000 11336 20052
rect 11388 20040 11394 20052
rect 13170 20040 13176 20052
rect 11388 20012 13176 20040
rect 11388 20000 11394 20012
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 13906 20000 13912 20052
rect 13964 20040 13970 20052
rect 14458 20040 14464 20052
rect 13964 20012 14464 20040
rect 13964 20000 13970 20012
rect 14458 20000 14464 20012
rect 14516 20040 14522 20052
rect 14826 20040 14832 20052
rect 14516 20012 14832 20040
rect 14516 20000 14522 20012
rect 14826 20000 14832 20012
rect 14884 20000 14890 20052
rect 22094 20040 22100 20052
rect 18524 20012 22100 20040
rect 4154 19932 4160 19984
rect 4212 19972 4218 19984
rect 14550 19972 14556 19984
rect 4212 19944 14556 19972
rect 4212 19932 4218 19944
rect 14550 19932 14556 19944
rect 14608 19932 14614 19984
rect 5626 19864 5632 19916
rect 5684 19904 5690 19916
rect 5813 19907 5871 19913
rect 5813 19904 5825 19907
rect 5684 19876 5825 19904
rect 5684 19864 5690 19876
rect 5813 19873 5825 19876
rect 5859 19873 5871 19907
rect 5813 19867 5871 19873
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19904 13783 19907
rect 14458 19904 14464 19916
rect 13771 19876 14464 19904
rect 13771 19873 13783 19876
rect 13725 19867 13783 19873
rect 14458 19864 14464 19876
rect 14516 19864 14522 19916
rect 18524 19913 18552 20012
rect 22094 20000 22100 20012
rect 22152 20000 22158 20052
rect 22186 20000 22192 20052
rect 22244 20040 22250 20052
rect 26326 20040 26332 20052
rect 22244 20012 26332 20040
rect 22244 20000 22250 20012
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 33042 20000 33048 20052
rect 33100 20000 33106 20052
rect 19306 19944 19564 19972
rect 18509 19907 18567 19913
rect 18509 19873 18521 19907
rect 18555 19873 18567 19907
rect 19306 19904 19334 19944
rect 18509 19867 18567 19873
rect 18616 19876 19334 19904
rect 19536 19904 19564 19944
rect 20346 19932 20352 19984
rect 20404 19972 20410 19984
rect 20404 19944 21036 19972
rect 20404 19932 20410 19944
rect 21008 19913 21036 19944
rect 21174 19932 21180 19984
rect 21232 19972 21238 19984
rect 21232 19944 22784 19972
rect 21232 19932 21238 19944
rect 20993 19907 21051 19913
rect 19536 19876 20668 19904
rect 2682 19796 2688 19848
rect 2740 19796 2746 19848
rect 5997 19839 6055 19845
rect 5997 19805 6009 19839
rect 6043 19836 6055 19839
rect 6178 19836 6184 19848
rect 6043 19808 6184 19836
rect 6043 19805 6055 19808
rect 5997 19799 6055 19805
rect 6178 19796 6184 19808
rect 6236 19796 6242 19848
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11606 19836 11612 19848
rect 11296 19808 11612 19836
rect 11296 19796 11302 19808
rect 11606 19796 11612 19808
rect 11664 19836 11670 19848
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 11664 19808 12449 19836
rect 11664 19796 11670 19808
rect 12437 19805 12449 19808
rect 12483 19836 12495 19839
rect 12526 19836 12532 19848
rect 12483 19808 12532 19836
rect 12483 19805 12495 19808
rect 12437 19799 12495 19805
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 12805 19839 12863 19845
rect 12805 19805 12817 19839
rect 12851 19836 12863 19839
rect 12894 19836 12900 19848
rect 12851 19808 12900 19836
rect 12851 19805 12863 19808
rect 12805 19799 12863 19805
rect 12894 19796 12900 19808
rect 12952 19796 12958 19848
rect 13173 19839 13231 19845
rect 13173 19805 13185 19839
rect 13219 19836 13231 19839
rect 13262 19836 13268 19848
rect 13219 19808 13268 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 13262 19796 13268 19808
rect 13320 19836 13326 19848
rect 17678 19836 17684 19848
rect 13320 19808 17684 19836
rect 13320 19796 13326 19808
rect 17678 19796 17684 19808
rect 17736 19836 17742 19848
rect 18616 19836 18644 19876
rect 17736 19808 18644 19836
rect 17736 19796 17742 19808
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 19288 19836 19294 19848
rect 18748 19808 19294 19836
rect 18748 19796 18754 19808
rect 19288 19796 19294 19808
rect 19346 19796 19352 19848
rect 20640 19845 20668 19876
rect 20993 19873 21005 19907
rect 21039 19873 21051 19907
rect 20993 19867 21051 19873
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 21726 19904 21732 19916
rect 21131 19876 21732 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 21726 19864 21732 19876
rect 21784 19864 21790 19916
rect 22370 19904 22376 19916
rect 21836 19876 22376 19904
rect 19439 19839 19497 19845
rect 19439 19805 19451 19839
rect 19485 19805 19497 19839
rect 19439 19799 19497 19805
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 20625 19839 20683 19845
rect 20625 19805 20637 19839
rect 20671 19836 20683 19839
rect 20714 19836 20720 19848
rect 20671 19808 20720 19836
rect 20671 19805 20683 19808
rect 20625 19799 20683 19805
rect 5445 19771 5503 19777
rect 5445 19737 5457 19771
rect 5491 19768 5503 19771
rect 5721 19771 5779 19777
rect 5721 19768 5733 19771
rect 5491 19740 5733 19768
rect 5491 19737 5503 19740
rect 5445 19731 5503 19737
rect 5721 19737 5733 19740
rect 5767 19768 5779 19771
rect 13630 19768 13636 19780
rect 5767 19740 13636 19768
rect 5767 19737 5779 19740
rect 5721 19731 5779 19737
rect 13630 19728 13636 19740
rect 13688 19728 13694 19780
rect 14369 19771 14427 19777
rect 14369 19737 14381 19771
rect 14415 19768 14427 19771
rect 17770 19768 17776 19780
rect 14415 19740 17776 19768
rect 14415 19737 14427 19740
rect 14369 19731 14427 19737
rect 17770 19728 17776 19740
rect 17828 19768 17834 19780
rect 19454 19768 19482 19799
rect 17828 19740 19482 19768
rect 17828 19728 17834 19740
rect 2777 19703 2835 19709
rect 2777 19669 2789 19703
rect 2823 19700 2835 19703
rect 4246 19700 4252 19712
rect 2823 19672 4252 19700
rect 2823 19669 2835 19672
rect 2777 19663 2835 19669
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 4430 19660 4436 19712
rect 4488 19700 4494 19712
rect 6181 19703 6239 19709
rect 6181 19700 6193 19703
rect 4488 19672 6193 19700
rect 4488 19660 4494 19672
rect 6181 19669 6193 19672
rect 6227 19669 6239 19703
rect 6181 19663 6239 19669
rect 12802 19660 12808 19712
rect 12860 19700 12866 19712
rect 14274 19700 14280 19712
rect 12860 19672 14280 19700
rect 12860 19660 12866 19672
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 14918 19660 14924 19712
rect 14976 19700 14982 19712
rect 17494 19700 17500 19712
rect 14976 19672 17500 19700
rect 14976 19660 14982 19672
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 18877 19703 18935 19709
rect 18877 19669 18889 19703
rect 18923 19700 18935 19703
rect 19242 19700 19248 19712
rect 18923 19672 19248 19700
rect 18923 19669 18935 19672
rect 18877 19663 18935 19669
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 19518 19660 19524 19712
rect 19576 19700 19582 19712
rect 19720 19700 19748 19799
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 21634 19796 21640 19848
rect 21692 19796 21698 19848
rect 21836 19845 21864 19876
rect 22370 19864 22376 19876
rect 22428 19864 22434 19916
rect 21821 19839 21879 19845
rect 21821 19805 21833 19839
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 22002 19796 22008 19848
rect 22060 19796 22066 19848
rect 22649 19839 22707 19845
rect 22649 19805 22661 19839
rect 22695 19834 22707 19839
rect 22756 19834 22784 19944
rect 22830 19932 22836 19984
rect 22888 19932 22894 19984
rect 31662 19904 31668 19916
rect 31312 19876 31668 19904
rect 22695 19806 22784 19834
rect 22695 19805 22707 19806
rect 22649 19799 22707 19805
rect 31018 19796 31024 19848
rect 31076 19836 31082 19848
rect 31312 19845 31340 19876
rect 31662 19864 31668 19876
rect 31720 19864 31726 19916
rect 31297 19839 31355 19845
rect 31297 19836 31309 19839
rect 31076 19808 31309 19836
rect 31076 19796 31082 19808
rect 31297 19805 31309 19808
rect 31343 19805 31355 19839
rect 31297 19799 31355 19805
rect 19794 19728 19800 19780
rect 19852 19768 19858 19780
rect 20533 19771 20591 19777
rect 20533 19768 20545 19771
rect 19852 19740 20545 19768
rect 19852 19728 19858 19740
rect 20533 19737 20545 19740
rect 20579 19737 20591 19771
rect 21913 19771 21971 19777
rect 21913 19768 21925 19771
rect 20533 19731 20591 19737
rect 21836 19740 21925 19768
rect 21836 19712 21864 19740
rect 21913 19737 21925 19740
rect 21959 19737 21971 19771
rect 21913 19731 21971 19737
rect 31573 19771 31631 19777
rect 31573 19737 31585 19771
rect 31619 19768 31631 19771
rect 31846 19768 31852 19780
rect 31619 19740 31852 19768
rect 31619 19737 31631 19740
rect 31573 19731 31631 19737
rect 31846 19728 31852 19740
rect 31904 19728 31910 19780
rect 32030 19728 32036 19780
rect 32088 19728 32094 19780
rect 19576 19672 19748 19700
rect 19576 19660 19582 19672
rect 21818 19660 21824 19712
rect 21876 19660 21882 19712
rect 22186 19660 22192 19712
rect 22244 19660 22250 19712
rect 25590 19660 25596 19712
rect 25648 19700 25654 19712
rect 36446 19700 36452 19712
rect 25648 19672 36452 19700
rect 25648 19660 25654 19672
rect 36446 19660 36452 19672
rect 36504 19660 36510 19712
rect 1104 19610 39352 19632
rect 1104 19558 10472 19610
rect 10524 19558 10536 19610
rect 10588 19558 10600 19610
rect 10652 19558 10664 19610
rect 10716 19558 10728 19610
rect 10780 19558 19994 19610
rect 20046 19558 20058 19610
rect 20110 19558 20122 19610
rect 20174 19558 20186 19610
rect 20238 19558 20250 19610
rect 20302 19558 29516 19610
rect 29568 19558 29580 19610
rect 29632 19558 29644 19610
rect 29696 19558 29708 19610
rect 29760 19558 29772 19610
rect 29824 19558 39038 19610
rect 39090 19558 39102 19610
rect 39154 19558 39166 19610
rect 39218 19558 39230 19610
rect 39282 19558 39294 19610
rect 39346 19558 39352 19610
rect 1104 19536 39352 19558
rect 9582 19496 9588 19508
rect 5460 19468 9588 19496
rect 3878 19388 3884 19440
rect 3936 19428 3942 19440
rect 4433 19431 4491 19437
rect 4433 19428 4445 19431
rect 3936 19400 4445 19428
rect 3936 19388 3942 19400
rect 4433 19397 4445 19400
rect 4479 19397 4491 19431
rect 4433 19391 4491 19397
rect 2682 19320 2688 19372
rect 2740 19360 2746 19372
rect 5460 19369 5488 19468
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 13998 19496 14004 19508
rect 13780 19468 14004 19496
rect 13780 19456 13786 19468
rect 13998 19456 14004 19468
rect 14056 19496 14062 19508
rect 14056 19468 14228 19496
rect 14056 19456 14062 19468
rect 5629 19431 5687 19437
rect 5629 19397 5641 19431
rect 5675 19428 5687 19431
rect 12986 19428 12992 19440
rect 5675 19400 12992 19428
rect 5675 19397 5687 19400
rect 5629 19391 5687 19397
rect 12986 19388 12992 19400
rect 13044 19388 13050 19440
rect 4341 19363 4399 19369
rect 4341 19360 4353 19363
rect 2740 19332 4353 19360
rect 2740 19320 2746 19332
rect 4341 19329 4353 19332
rect 4387 19360 4399 19363
rect 5445 19363 5503 19369
rect 4387 19332 5396 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 5368 19292 5396 19332
rect 5445 19329 5457 19363
rect 5491 19329 5503 19363
rect 5445 19323 5503 19329
rect 5721 19363 5779 19369
rect 5721 19329 5733 19363
rect 5767 19329 5779 19363
rect 5721 19323 5779 19329
rect 5813 19363 5871 19369
rect 5813 19329 5825 19363
rect 5859 19360 5871 19363
rect 11330 19360 11336 19372
rect 5859 19332 11336 19360
rect 5859 19329 5871 19332
rect 5813 19323 5871 19329
rect 5626 19292 5632 19304
rect 5368 19264 5632 19292
rect 5626 19252 5632 19264
rect 5684 19252 5690 19304
rect 5166 19184 5172 19236
rect 5224 19224 5230 19236
rect 5736 19224 5764 19323
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19360 11943 19363
rect 12250 19360 12256 19372
rect 11931 19332 12256 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 12250 19320 12256 19332
rect 12308 19320 12314 19372
rect 12434 19320 12440 19372
rect 12492 19320 12498 19372
rect 13814 19320 13820 19372
rect 13872 19320 13878 19372
rect 14200 19360 14228 19468
rect 14274 19456 14280 19508
rect 14332 19496 14338 19508
rect 15289 19499 15347 19505
rect 14332 19468 15056 19496
rect 14332 19456 14338 19468
rect 14918 19388 14924 19440
rect 14976 19388 14982 19440
rect 15028 19437 15056 19468
rect 15289 19465 15301 19499
rect 15335 19496 15347 19499
rect 20099 19499 20157 19505
rect 15335 19468 20024 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 15013 19431 15071 19437
rect 15013 19397 15025 19431
rect 15059 19397 15071 19431
rect 15013 19391 15071 19397
rect 16666 19388 16672 19440
rect 16724 19428 16730 19440
rect 19794 19428 19800 19440
rect 16724 19400 19800 19428
rect 16724 19388 16730 19400
rect 19794 19388 19800 19400
rect 19852 19388 19858 19440
rect 19886 19388 19892 19440
rect 19944 19388 19950 19440
rect 19996 19428 20024 19468
rect 20099 19465 20111 19499
rect 20145 19496 20157 19499
rect 21082 19496 21088 19508
rect 20145 19468 21088 19496
rect 20145 19465 20157 19468
rect 20099 19459 20157 19465
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 21726 19456 21732 19508
rect 21784 19496 21790 19508
rect 22002 19496 22008 19508
rect 21784 19468 22008 19496
rect 21784 19456 21790 19468
rect 22002 19456 22008 19468
rect 22060 19456 22066 19508
rect 24578 19496 24584 19508
rect 22388 19468 24584 19496
rect 20438 19428 20444 19440
rect 19996 19400 20444 19428
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 14200 19332 14749 19360
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 15105 19363 15163 19369
rect 15105 19360 15117 19363
rect 14884 19332 15117 19360
rect 14884 19320 14890 19332
rect 15105 19329 15117 19332
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 17218 19320 17224 19372
rect 17276 19360 17282 19372
rect 17497 19363 17555 19369
rect 17497 19360 17509 19363
rect 17276 19332 17509 19360
rect 17276 19320 17282 19332
rect 17497 19329 17509 19332
rect 17543 19329 17555 19363
rect 17497 19323 17555 19329
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19360 17647 19363
rect 18138 19360 18144 19372
rect 17635 19332 18144 19360
rect 17635 19329 17647 19332
rect 17589 19323 17647 19329
rect 18138 19320 18144 19332
rect 18196 19320 18202 19372
rect 18782 19320 18788 19372
rect 18840 19360 18846 19372
rect 18966 19360 18972 19372
rect 18840 19332 18972 19360
rect 18840 19320 18846 19332
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 20530 19360 20536 19372
rect 19484 19332 20536 19360
rect 19484 19320 19490 19332
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 20772 19332 20821 19360
rect 20772 19320 20778 19332
rect 20809 19329 20821 19332
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 22278 19320 22284 19372
rect 22336 19360 22342 19372
rect 22388 19369 22416 19468
rect 24578 19456 24584 19468
rect 24636 19456 24642 19508
rect 24762 19456 24768 19508
rect 24820 19496 24826 19508
rect 26329 19499 26387 19505
rect 26329 19496 26341 19499
rect 24820 19468 26341 19496
rect 24820 19456 24826 19468
rect 26329 19465 26341 19468
rect 26375 19496 26387 19499
rect 27522 19496 27528 19508
rect 26375 19468 27528 19496
rect 26375 19465 26387 19468
rect 26329 19459 26387 19465
rect 27522 19456 27528 19468
rect 27580 19456 27586 19508
rect 28166 19456 28172 19508
rect 28224 19496 28230 19508
rect 31297 19499 31355 19505
rect 28224 19468 31064 19496
rect 28224 19456 28230 19468
rect 23934 19428 23940 19440
rect 23874 19400 23940 19428
rect 23934 19388 23940 19400
rect 23992 19388 23998 19440
rect 30650 19428 30656 19440
rect 26082 19400 30656 19428
rect 30650 19388 30656 19400
rect 30708 19388 30714 19440
rect 31036 19437 31064 19468
rect 31297 19465 31309 19499
rect 31343 19496 31355 19499
rect 31343 19468 32996 19496
rect 31343 19465 31355 19468
rect 31297 19459 31355 19465
rect 31021 19431 31079 19437
rect 31021 19397 31033 19431
rect 31067 19397 31079 19431
rect 32968 19428 32996 19468
rect 33134 19456 33140 19508
rect 33192 19496 33198 19508
rect 36081 19499 36139 19505
rect 36081 19496 36093 19499
rect 33192 19468 36093 19496
rect 33192 19456 33198 19468
rect 36081 19465 36093 19468
rect 36127 19465 36139 19499
rect 36081 19459 36139 19465
rect 36446 19456 36452 19508
rect 36504 19456 36510 19508
rect 33226 19428 33232 19440
rect 32968 19400 33232 19428
rect 31021 19391 31079 19397
rect 33226 19388 33232 19400
rect 33284 19388 33290 19440
rect 33778 19388 33784 19440
rect 33836 19428 33842 19440
rect 35437 19431 35495 19437
rect 35437 19428 35449 19431
rect 33836 19400 35449 19428
rect 33836 19388 33842 19400
rect 35437 19397 35449 19400
rect 35483 19397 35495 19431
rect 35437 19391 35495 19397
rect 35529 19431 35587 19437
rect 35529 19397 35541 19431
rect 35575 19428 35587 19431
rect 35894 19428 35900 19440
rect 35575 19400 35900 19428
rect 35575 19397 35587 19400
rect 35529 19391 35587 19397
rect 35894 19388 35900 19400
rect 35952 19388 35958 19440
rect 22373 19363 22431 19369
rect 22373 19360 22385 19363
rect 22336 19332 22385 19360
rect 22336 19320 22342 19332
rect 22373 19329 22385 19332
rect 22419 19329 22431 19363
rect 22373 19323 22431 19329
rect 24578 19320 24584 19372
rect 24636 19320 24642 19372
rect 30742 19320 30748 19372
rect 30800 19320 30806 19372
rect 30834 19320 30840 19372
rect 30892 19360 30898 19372
rect 30929 19363 30987 19369
rect 30929 19360 30941 19363
rect 30892 19332 30941 19360
rect 30892 19320 30898 19332
rect 30929 19329 30941 19332
rect 30975 19329 30987 19363
rect 30929 19323 30987 19329
rect 31110 19320 31116 19372
rect 31168 19320 31174 19372
rect 34974 19320 34980 19372
rect 35032 19360 35038 19372
rect 35253 19363 35311 19369
rect 35253 19360 35265 19363
rect 35032 19332 35265 19360
rect 35032 19320 35038 19332
rect 35253 19329 35265 19332
rect 35299 19329 35311 19363
rect 35253 19323 35311 19329
rect 35618 19320 35624 19372
rect 35676 19360 35682 19372
rect 36541 19363 36599 19369
rect 36541 19360 36553 19363
rect 35676 19332 36553 19360
rect 35676 19320 35682 19332
rect 36541 19329 36553 19332
rect 36587 19329 36599 19363
rect 36541 19323 36599 19329
rect 12710 19252 12716 19304
rect 12768 19252 12774 19304
rect 21174 19292 21180 19304
rect 17236 19264 21180 19292
rect 5224 19196 5764 19224
rect 5224 19184 5230 19196
rect 5994 19184 6000 19236
rect 6052 19184 6058 19236
rect 14185 19227 14243 19233
rect 14185 19193 14197 19227
rect 14231 19224 14243 19227
rect 14274 19224 14280 19236
rect 14231 19196 14280 19224
rect 14231 19193 14243 19196
rect 14185 19187 14243 19193
rect 14274 19184 14280 19196
rect 14332 19184 14338 19236
rect 2222 19116 2228 19168
rect 2280 19156 2286 19168
rect 6086 19156 6092 19168
rect 2280 19128 6092 19156
rect 2280 19116 2286 19128
rect 6086 19116 6092 19128
rect 6144 19116 6150 19168
rect 11885 19159 11943 19165
rect 11885 19125 11897 19159
rect 11931 19156 11943 19159
rect 17236 19156 17264 19264
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 21358 19252 21364 19304
rect 21416 19252 21422 19304
rect 22646 19252 22652 19304
rect 22704 19252 22710 19304
rect 24857 19295 24915 19301
rect 24857 19261 24869 19295
rect 24903 19292 24915 19295
rect 27154 19292 27160 19304
rect 24903 19264 27160 19292
rect 24903 19261 24915 19264
rect 24857 19255 24915 19261
rect 27154 19252 27160 19264
rect 27212 19252 27218 19304
rect 27890 19252 27896 19304
rect 27948 19292 27954 19304
rect 28534 19292 28540 19304
rect 27948 19264 28540 19292
rect 27948 19252 27954 19264
rect 28534 19252 28540 19264
rect 28592 19292 28598 19304
rect 36633 19295 36691 19301
rect 28592 19264 31754 19292
rect 28592 19252 28598 19264
rect 22094 19224 22100 19236
rect 20088 19196 22100 19224
rect 20088 19165 20116 19196
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 31726 19224 31754 19264
rect 36633 19261 36645 19295
rect 36679 19261 36691 19295
rect 36633 19255 36691 19261
rect 36648 19224 36676 19255
rect 37458 19224 37464 19236
rect 23676 19196 24256 19224
rect 11931 19128 17264 19156
rect 20073 19159 20131 19165
rect 11931 19125 11943 19128
rect 11885 19119 11943 19125
rect 20073 19125 20085 19159
rect 20119 19125 20131 19159
rect 20073 19119 20131 19125
rect 20257 19159 20315 19165
rect 20257 19125 20269 19159
rect 20303 19156 20315 19159
rect 20530 19156 20536 19168
rect 20303 19128 20536 19156
rect 20303 19125 20315 19128
rect 20257 19119 20315 19125
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 23676 19156 23704 19196
rect 21232 19128 23704 19156
rect 21232 19116 21238 19128
rect 24118 19116 24124 19168
rect 24176 19116 24182 19168
rect 24228 19156 24256 19196
rect 28966 19196 31432 19224
rect 31726 19196 37464 19224
rect 28966 19156 28994 19196
rect 24228 19128 28994 19156
rect 31404 19156 31432 19196
rect 37458 19184 37464 19196
rect 37516 19184 37522 19236
rect 34606 19156 34612 19168
rect 31404 19128 34612 19156
rect 34606 19116 34612 19128
rect 34664 19116 34670 19168
rect 34698 19116 34704 19168
rect 34756 19156 34762 19168
rect 34977 19159 35035 19165
rect 34977 19156 34989 19159
rect 34756 19128 34989 19156
rect 34756 19116 34762 19128
rect 34977 19125 34989 19128
rect 35023 19125 35035 19159
rect 34977 19119 35035 19125
rect 1104 19066 39192 19088
rect 1104 19014 5711 19066
rect 5763 19014 5775 19066
rect 5827 19014 5839 19066
rect 5891 19014 5903 19066
rect 5955 19014 5967 19066
rect 6019 19014 15233 19066
rect 15285 19014 15297 19066
rect 15349 19014 15361 19066
rect 15413 19014 15425 19066
rect 15477 19014 15489 19066
rect 15541 19014 24755 19066
rect 24807 19014 24819 19066
rect 24871 19014 24883 19066
rect 24935 19014 24947 19066
rect 24999 19014 25011 19066
rect 25063 19014 34277 19066
rect 34329 19014 34341 19066
rect 34393 19014 34405 19066
rect 34457 19014 34469 19066
rect 34521 19014 34533 19066
rect 34585 19014 39192 19066
rect 1104 18992 39192 19014
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21726 18952 21732 18964
rect 20772 18924 21732 18952
rect 20772 18912 20778 18924
rect 21726 18912 21732 18924
rect 21784 18952 21790 18964
rect 26602 18952 26608 18964
rect 21784 18924 26608 18952
rect 21784 18912 21790 18924
rect 26602 18912 26608 18924
rect 26660 18912 26666 18964
rect 27798 18912 27804 18964
rect 27856 18952 27862 18964
rect 28261 18955 28319 18961
rect 28261 18952 28273 18955
rect 27856 18924 28273 18952
rect 27856 18912 27862 18924
rect 28261 18921 28273 18924
rect 28307 18921 28319 18955
rect 35434 18952 35440 18964
rect 28261 18915 28319 18921
rect 28368 18924 35440 18952
rect 25498 18844 25504 18896
rect 25556 18884 25562 18896
rect 25556 18856 26556 18884
rect 25556 18844 25562 18856
rect 20809 18819 20867 18825
rect 20809 18785 20821 18819
rect 20855 18816 20867 18819
rect 22278 18816 22284 18828
rect 20855 18788 22284 18816
rect 20855 18785 20867 18788
rect 20809 18779 20867 18785
rect 22278 18776 22284 18788
rect 22336 18776 22342 18828
rect 23661 18819 23719 18825
rect 23661 18785 23673 18819
rect 23707 18816 23719 18819
rect 25130 18816 25136 18828
rect 23707 18788 25136 18816
rect 23707 18785 23719 18788
rect 23661 18779 23719 18785
rect 25130 18776 25136 18788
rect 25188 18776 25194 18828
rect 25406 18776 25412 18828
rect 25464 18816 25470 18828
rect 26237 18819 26295 18825
rect 26237 18816 26249 18819
rect 25464 18788 26249 18816
rect 25464 18776 25470 18788
rect 26237 18785 26249 18788
rect 26283 18785 26295 18819
rect 26237 18779 26295 18785
rect 26326 18776 26332 18828
rect 26384 18776 26390 18828
rect 26418 18776 26424 18828
rect 26476 18776 26482 18828
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 4430 18748 4436 18760
rect 1719 18720 4436 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 4430 18708 4436 18720
rect 4488 18708 4494 18760
rect 5626 18708 5632 18760
rect 5684 18748 5690 18760
rect 6273 18751 6331 18757
rect 6273 18748 6285 18751
rect 5684 18720 6285 18748
rect 5684 18708 5690 18720
rect 6273 18717 6285 18720
rect 6319 18748 6331 18751
rect 6546 18748 6552 18760
rect 6319 18720 6552 18748
rect 6319 18717 6331 18720
rect 6273 18711 6331 18717
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12250 18748 12256 18760
rect 12115 18720 12256 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 19702 18708 19708 18760
rect 19760 18748 19766 18760
rect 19889 18751 19947 18757
rect 19889 18748 19901 18751
rect 19760 18720 19901 18748
rect 19760 18708 19766 18720
rect 19889 18717 19901 18720
rect 19935 18717 19947 18751
rect 19889 18711 19947 18717
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 23477 18751 23535 18757
rect 23477 18748 23489 18751
rect 22796 18720 23489 18748
rect 22796 18708 22802 18720
rect 23477 18717 23489 18720
rect 23523 18717 23535 18751
rect 23477 18711 23535 18717
rect 24949 18751 25007 18757
rect 24949 18717 24961 18751
rect 24995 18748 25007 18751
rect 26528 18748 26556 18856
rect 27062 18844 27068 18896
rect 27120 18844 27126 18896
rect 28368 18884 28396 18924
rect 35434 18912 35440 18924
rect 35492 18952 35498 18964
rect 35492 18924 35940 18952
rect 35492 18912 35498 18924
rect 27172 18856 28396 18884
rect 26786 18776 26792 18828
rect 26844 18816 26850 18828
rect 27172 18816 27200 18856
rect 30650 18844 30656 18896
rect 30708 18844 30714 18896
rect 26844 18788 27200 18816
rect 27525 18819 27583 18825
rect 26844 18776 26850 18788
rect 27525 18785 27537 18819
rect 27571 18816 27583 18819
rect 30466 18816 30472 18828
rect 27571 18788 30472 18816
rect 27571 18785 27583 18788
rect 27525 18779 27583 18785
rect 30466 18776 30472 18788
rect 30524 18776 30530 18828
rect 31018 18776 31024 18828
rect 31076 18816 31082 18828
rect 32309 18819 32367 18825
rect 32309 18816 32321 18819
rect 31076 18788 32321 18816
rect 31076 18776 31082 18788
rect 32309 18785 32321 18788
rect 32355 18785 32367 18819
rect 32309 18779 32367 18785
rect 32585 18819 32643 18825
rect 32585 18785 32597 18819
rect 32631 18816 32643 18819
rect 33134 18816 33140 18828
rect 32631 18788 33140 18816
rect 32631 18785 32643 18788
rect 32585 18779 32643 18785
rect 33134 18776 33140 18788
rect 33192 18776 33198 18828
rect 34333 18819 34391 18825
rect 34333 18785 34345 18819
rect 34379 18816 34391 18819
rect 35618 18816 35624 18828
rect 34379 18788 35624 18816
rect 34379 18785 34391 18788
rect 34333 18779 34391 18785
rect 28169 18751 28227 18757
rect 28169 18748 28181 18751
rect 24995 18720 26464 18748
rect 26528 18720 28181 18748
rect 24995 18717 25007 18720
rect 24949 18711 25007 18717
rect 2866 18640 2872 18692
rect 2924 18680 2930 18692
rect 6365 18683 6423 18689
rect 6365 18680 6377 18683
rect 2924 18652 6377 18680
rect 2924 18640 2930 18652
rect 6365 18649 6377 18652
rect 6411 18649 6423 18683
rect 6365 18643 6423 18649
rect 17770 18640 17776 18692
rect 17828 18640 17834 18692
rect 17862 18640 17868 18692
rect 17920 18680 17926 18692
rect 18509 18683 18567 18689
rect 18509 18680 18521 18683
rect 17920 18652 18521 18680
rect 17920 18640 17926 18652
rect 18509 18649 18521 18652
rect 18555 18649 18567 18683
rect 18509 18643 18567 18649
rect 19518 18640 19524 18692
rect 19576 18680 19582 18692
rect 20165 18683 20223 18689
rect 20165 18680 20177 18683
rect 19576 18652 20177 18680
rect 19576 18640 19582 18652
rect 20165 18649 20177 18652
rect 20211 18649 20223 18683
rect 20165 18643 20223 18649
rect 21082 18640 21088 18692
rect 21140 18640 21146 18692
rect 24026 18680 24032 18692
rect 22310 18652 24032 18680
rect 24026 18640 24032 18652
rect 24084 18640 24090 18692
rect 25406 18640 25412 18692
rect 25464 18640 25470 18692
rect 26436 18680 26464 18720
rect 28169 18717 28181 18720
rect 28215 18717 28227 18751
rect 28169 18711 28227 18717
rect 28258 18708 28264 18760
rect 28316 18748 28322 18760
rect 28316 18720 31754 18748
rect 28316 18708 28322 18720
rect 26878 18680 26884 18692
rect 26436 18652 26884 18680
rect 26878 18640 26884 18652
rect 26936 18640 26942 18692
rect 27617 18683 27675 18689
rect 27617 18649 27629 18683
rect 27663 18680 27675 18683
rect 27890 18680 27896 18692
rect 27663 18652 27896 18680
rect 27663 18649 27675 18652
rect 27617 18643 27675 18649
rect 27890 18640 27896 18652
rect 27948 18640 27954 18692
rect 30834 18640 30840 18692
rect 30892 18680 30898 18692
rect 30929 18683 30987 18689
rect 30929 18680 30941 18683
rect 30892 18652 30941 18680
rect 30892 18640 30898 18652
rect 30929 18649 30941 18652
rect 30975 18649 30987 18683
rect 30929 18643 30987 18649
rect 31202 18640 31208 18692
rect 31260 18640 31266 18692
rect 934 18572 940 18624
rect 992 18612 998 18624
rect 1765 18615 1823 18621
rect 1765 18612 1777 18615
rect 992 18584 1777 18612
rect 992 18572 998 18584
rect 1765 18581 1777 18584
rect 1811 18581 1823 18615
rect 1765 18575 1823 18581
rect 5718 18572 5724 18624
rect 5776 18572 5782 18624
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 12161 18615 12219 18621
rect 12161 18612 12173 18615
rect 9088 18584 12173 18612
rect 9088 18572 9094 18584
rect 12161 18581 12173 18584
rect 12207 18581 12219 18615
rect 12161 18575 12219 18581
rect 21726 18572 21732 18624
rect 21784 18612 21790 18624
rect 22557 18615 22615 18621
rect 22557 18612 22569 18615
rect 21784 18584 22569 18612
rect 21784 18572 21790 18584
rect 22557 18581 22569 18584
rect 22603 18581 22615 18615
rect 22557 18575 22615 18581
rect 23014 18572 23020 18624
rect 23072 18572 23078 18624
rect 23382 18572 23388 18624
rect 23440 18572 23446 18624
rect 26053 18615 26111 18621
rect 26053 18581 26065 18615
rect 26099 18612 26111 18615
rect 27154 18612 27160 18624
rect 26099 18584 27160 18612
rect 26099 18581 26111 18584
rect 26053 18575 26111 18581
rect 27154 18572 27160 18584
rect 27212 18572 27218 18624
rect 27522 18572 27528 18624
rect 27580 18572 27586 18624
rect 30742 18572 30748 18624
rect 30800 18612 30806 18624
rect 31113 18615 31171 18621
rect 31113 18612 31125 18615
rect 30800 18584 31125 18612
rect 30800 18572 30806 18584
rect 31113 18581 31125 18584
rect 31159 18612 31171 18615
rect 31294 18612 31300 18624
rect 31159 18584 31300 18612
rect 31159 18581 31171 18584
rect 31113 18575 31171 18581
rect 31294 18572 31300 18584
rect 31352 18572 31358 18624
rect 31726 18612 31754 18720
rect 34054 18680 34060 18692
rect 33810 18652 34060 18680
rect 34054 18640 34060 18652
rect 34112 18640 34118 18692
rect 34348 18612 34376 18779
rect 35618 18776 35624 18788
rect 35676 18776 35682 18828
rect 35710 18708 35716 18760
rect 35768 18708 35774 18760
rect 35912 18748 35940 18924
rect 37458 18776 37464 18828
rect 37516 18776 37522 18828
rect 37185 18751 37243 18757
rect 37185 18748 37197 18751
rect 35912 18720 37197 18748
rect 37185 18717 37197 18720
rect 37231 18717 37243 18751
rect 37185 18711 37243 18717
rect 36449 18683 36507 18689
rect 36449 18649 36461 18683
rect 36495 18680 36507 18683
rect 36814 18680 36820 18692
rect 36495 18652 36820 18680
rect 36495 18649 36507 18652
rect 36449 18643 36507 18649
rect 36814 18640 36820 18652
rect 36872 18640 36878 18692
rect 31726 18584 34376 18612
rect 1104 18522 39352 18544
rect 1104 18470 10472 18522
rect 10524 18470 10536 18522
rect 10588 18470 10600 18522
rect 10652 18470 10664 18522
rect 10716 18470 10728 18522
rect 10780 18470 19994 18522
rect 20046 18470 20058 18522
rect 20110 18470 20122 18522
rect 20174 18470 20186 18522
rect 20238 18470 20250 18522
rect 20302 18470 29516 18522
rect 29568 18470 29580 18522
rect 29632 18470 29644 18522
rect 29696 18470 29708 18522
rect 29760 18470 29772 18522
rect 29824 18470 39038 18522
rect 39090 18470 39102 18522
rect 39154 18470 39166 18522
rect 39218 18470 39230 18522
rect 39282 18470 39294 18522
rect 39346 18470 39352 18522
rect 1104 18448 39352 18470
rect 5718 18368 5724 18420
rect 5776 18408 5782 18420
rect 17954 18408 17960 18420
rect 5776 18380 17264 18408
rect 5776 18368 5782 18380
rect 2958 18300 2964 18352
rect 3016 18300 3022 18352
rect 3694 18300 3700 18352
rect 3752 18300 3758 18352
rect 11238 18300 11244 18352
rect 11296 18340 11302 18352
rect 11296 18312 13938 18340
rect 11296 18300 11302 18312
rect 12434 18232 12440 18284
rect 12492 18272 12498 18284
rect 13170 18272 13176 18284
rect 12492 18244 13176 18272
rect 12492 18232 12498 18244
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2685 18207 2743 18213
rect 2685 18204 2697 18207
rect 2280 18176 2697 18204
rect 2280 18164 2286 18176
rect 2685 18173 2697 18176
rect 2731 18173 2743 18207
rect 2685 18167 2743 18173
rect 4433 18207 4491 18213
rect 4433 18173 4445 18207
rect 4479 18204 4491 18207
rect 6914 18204 6920 18216
rect 4479 18176 6920 18204
rect 4479 18173 4491 18176
rect 4433 18167 4491 18173
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 13449 18207 13507 18213
rect 13449 18173 13461 18207
rect 13495 18204 13507 18207
rect 14734 18204 14740 18216
rect 13495 18176 14740 18204
rect 13495 18173 13507 18176
rect 13449 18167 13507 18173
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 17236 18204 17264 18380
rect 17328 18380 17960 18408
rect 17328 18281 17356 18380
rect 17954 18368 17960 18380
rect 18012 18408 18018 18420
rect 19426 18408 19432 18420
rect 18012 18380 19432 18408
rect 18012 18368 18018 18380
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 20622 18368 20628 18420
rect 20680 18368 20686 18420
rect 21269 18411 21327 18417
rect 21269 18377 21281 18411
rect 21315 18408 21327 18411
rect 22738 18408 22744 18420
rect 21315 18380 22744 18408
rect 21315 18377 21327 18380
rect 21269 18371 21327 18377
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 24026 18368 24032 18420
rect 24084 18368 24090 18420
rect 24486 18368 24492 18420
rect 24544 18408 24550 18420
rect 24581 18411 24639 18417
rect 24581 18408 24593 18411
rect 24544 18380 24593 18408
rect 24544 18368 24550 18380
rect 24581 18377 24593 18380
rect 24627 18377 24639 18411
rect 24581 18371 24639 18377
rect 25041 18411 25099 18417
rect 25041 18377 25053 18411
rect 25087 18408 25099 18411
rect 26510 18408 26516 18420
rect 25087 18380 26516 18408
rect 25087 18377 25099 18380
rect 25041 18371 25099 18377
rect 26510 18368 26516 18380
rect 26568 18368 26574 18420
rect 30650 18368 30656 18420
rect 30708 18408 30714 18420
rect 31297 18411 31355 18417
rect 31297 18408 31309 18411
rect 30708 18380 31309 18408
rect 30708 18368 30714 18380
rect 31297 18377 31309 18380
rect 31343 18408 31355 18411
rect 32582 18408 32588 18420
rect 31343 18380 32588 18408
rect 31343 18377 31355 18380
rect 31297 18371 31355 18377
rect 32582 18368 32588 18380
rect 32640 18368 32646 18420
rect 37182 18368 37188 18420
rect 37240 18408 37246 18420
rect 37553 18411 37611 18417
rect 37553 18408 37565 18411
rect 37240 18380 37565 18408
rect 37240 18368 37246 18380
rect 37553 18377 37565 18380
rect 37599 18377 37611 18411
rect 37553 18371 37611 18377
rect 17494 18300 17500 18352
rect 17552 18300 17558 18352
rect 19518 18300 19524 18352
rect 19576 18340 19582 18352
rect 19797 18343 19855 18349
rect 19797 18340 19809 18343
rect 19576 18312 19809 18340
rect 19576 18300 19582 18312
rect 19797 18309 19809 18312
rect 19843 18309 19855 18343
rect 19797 18303 19855 18309
rect 19889 18343 19947 18349
rect 19889 18309 19901 18343
rect 19935 18340 19947 18343
rect 31205 18343 31263 18349
rect 31205 18340 31217 18343
rect 19935 18312 31217 18340
rect 19935 18309 19947 18312
rect 19889 18303 19947 18309
rect 31205 18309 31217 18312
rect 31251 18340 31263 18343
rect 31570 18340 31576 18352
rect 31251 18312 31576 18340
rect 31251 18309 31263 18312
rect 31205 18303 31263 18309
rect 31570 18300 31576 18312
rect 31628 18300 31634 18352
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18241 17371 18275
rect 17313 18235 17371 18241
rect 17586 18232 17592 18284
rect 17644 18232 17650 18284
rect 17681 18275 17739 18281
rect 17681 18241 17693 18275
rect 17727 18272 17739 18275
rect 17862 18272 17868 18284
rect 17727 18244 17868 18272
rect 17727 18241 17739 18244
rect 17681 18235 17739 18241
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 18874 18232 18880 18284
rect 18932 18272 18938 18284
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 18932 18244 19625 18272
rect 18932 18232 18938 18244
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 19978 18232 19984 18284
rect 20036 18232 20042 18284
rect 20530 18232 20536 18284
rect 20588 18272 20594 18284
rect 20901 18275 20959 18281
rect 20901 18272 20913 18275
rect 20588 18244 20913 18272
rect 20588 18232 20594 18244
rect 20901 18241 20913 18244
rect 20947 18241 20959 18275
rect 20901 18235 20959 18241
rect 21358 18232 21364 18284
rect 21416 18272 21422 18284
rect 22557 18275 22615 18281
rect 21416 18244 22094 18272
rect 21416 18232 21422 18244
rect 22066 18204 22094 18244
rect 22557 18241 22569 18275
rect 22603 18272 22615 18275
rect 22646 18272 22652 18284
rect 22603 18244 22652 18272
rect 22603 18241 22615 18244
rect 22557 18235 22615 18241
rect 22646 18232 22652 18244
rect 22704 18232 22710 18284
rect 22830 18232 22836 18284
rect 22888 18272 22894 18284
rect 22888 18244 23336 18272
rect 22888 18232 22894 18244
rect 23198 18204 23204 18216
rect 17236 18176 21220 18204
rect 22066 18176 23204 18204
rect 20165 18139 20223 18145
rect 20165 18105 20177 18139
rect 20211 18136 20223 18139
rect 21085 18139 21143 18145
rect 21085 18136 21097 18139
rect 20211 18108 21097 18136
rect 20211 18105 20223 18108
rect 20165 18099 20223 18105
rect 21085 18105 21097 18108
rect 21131 18105 21143 18139
rect 21192 18136 21220 18176
rect 23198 18164 23204 18176
rect 23256 18164 23262 18216
rect 23308 18213 23336 18244
rect 23382 18232 23388 18284
rect 23440 18272 23446 18284
rect 23937 18275 23995 18281
rect 23937 18272 23949 18275
rect 23440 18244 23949 18272
rect 23440 18232 23446 18244
rect 23937 18241 23949 18244
rect 23983 18241 23995 18275
rect 23937 18235 23995 18241
rect 24949 18275 25007 18281
rect 24949 18241 24961 18275
rect 24995 18272 25007 18275
rect 25314 18272 25320 18284
rect 24995 18244 25320 18272
rect 24995 18241 25007 18244
rect 24949 18235 25007 18241
rect 25314 18232 25320 18244
rect 25372 18232 25378 18284
rect 25866 18232 25872 18284
rect 25924 18232 25930 18284
rect 26602 18232 26608 18284
rect 26660 18232 26666 18284
rect 27154 18232 27160 18284
rect 27212 18232 27218 18284
rect 30834 18232 30840 18284
rect 30892 18272 30898 18284
rect 31478 18272 31484 18284
rect 30892 18244 31484 18272
rect 30892 18232 30898 18244
rect 31478 18232 31484 18244
rect 31536 18232 31542 18284
rect 33962 18232 33968 18284
rect 34020 18272 34026 18284
rect 35621 18275 35679 18281
rect 35621 18272 35633 18275
rect 34020 18244 35633 18272
rect 34020 18232 34026 18244
rect 35621 18241 35633 18244
rect 35667 18272 35679 18275
rect 36814 18272 36820 18284
rect 35667 18244 36820 18272
rect 35667 18241 35679 18244
rect 35621 18235 35679 18241
rect 36814 18232 36820 18244
rect 36872 18232 36878 18284
rect 37182 18232 37188 18284
rect 37240 18272 37246 18284
rect 37461 18275 37519 18281
rect 37461 18272 37473 18275
rect 37240 18244 37473 18272
rect 37240 18232 37246 18244
rect 37461 18241 37473 18244
rect 37507 18241 37519 18275
rect 37461 18235 37519 18241
rect 23293 18207 23351 18213
rect 23293 18173 23305 18207
rect 23339 18204 23351 18207
rect 23750 18204 23756 18216
rect 23339 18176 23756 18204
rect 23339 18173 23351 18176
rect 23293 18167 23351 18173
rect 23750 18164 23756 18176
rect 23808 18164 23814 18216
rect 25130 18164 25136 18216
rect 25188 18164 25194 18216
rect 26326 18164 26332 18216
rect 26384 18164 26390 18216
rect 26620 18204 26648 18232
rect 27341 18207 27399 18213
rect 27341 18204 27353 18207
rect 26620 18176 27353 18204
rect 27341 18173 27353 18176
rect 27387 18173 27399 18207
rect 27341 18167 27399 18173
rect 27706 18164 27712 18216
rect 27764 18204 27770 18216
rect 31202 18204 31208 18216
rect 27764 18176 31208 18204
rect 27764 18164 27770 18176
rect 31202 18164 31208 18176
rect 31260 18204 31266 18216
rect 31389 18207 31447 18213
rect 31389 18204 31401 18207
rect 31260 18176 31401 18204
rect 31260 18164 31266 18176
rect 31389 18173 31401 18176
rect 31435 18204 31447 18207
rect 34146 18204 34152 18216
rect 31435 18176 34152 18204
rect 31435 18173 31447 18176
rect 31389 18167 31447 18173
rect 34146 18164 34152 18176
rect 34204 18164 34210 18216
rect 35894 18164 35900 18216
rect 35952 18204 35958 18216
rect 36446 18204 36452 18216
rect 35952 18176 36452 18204
rect 35952 18164 35958 18176
rect 36446 18164 36452 18176
rect 36504 18164 36510 18216
rect 26050 18136 26056 18148
rect 21192 18108 26056 18136
rect 21085 18099 21143 18105
rect 26050 18096 26056 18108
rect 26108 18096 26114 18148
rect 14918 18028 14924 18080
rect 14976 18028 14982 18080
rect 17862 18028 17868 18080
rect 17920 18028 17926 18080
rect 20438 18028 20444 18080
rect 20496 18068 20502 18080
rect 20993 18071 21051 18077
rect 20993 18068 21005 18071
rect 20496 18040 21005 18068
rect 20496 18028 20502 18040
rect 20993 18037 21005 18040
rect 21039 18037 21051 18071
rect 20993 18031 21051 18037
rect 26142 18028 26148 18080
rect 26200 18028 26206 18080
rect 26237 18071 26295 18077
rect 26237 18037 26249 18071
rect 26283 18068 26295 18071
rect 26970 18068 26976 18080
rect 26283 18040 26976 18068
rect 26283 18037 26295 18040
rect 26237 18031 26295 18037
rect 26970 18028 26976 18040
rect 27028 18028 27034 18080
rect 30837 18071 30895 18077
rect 30837 18037 30849 18071
rect 30883 18068 30895 18071
rect 31294 18068 31300 18080
rect 30883 18040 31300 18068
rect 30883 18037 30895 18040
rect 30837 18031 30895 18037
rect 31294 18028 31300 18040
rect 31352 18028 31358 18080
rect 1104 17978 39192 18000
rect 1104 17926 5711 17978
rect 5763 17926 5775 17978
rect 5827 17926 5839 17978
rect 5891 17926 5903 17978
rect 5955 17926 5967 17978
rect 6019 17926 15233 17978
rect 15285 17926 15297 17978
rect 15349 17926 15361 17978
rect 15413 17926 15425 17978
rect 15477 17926 15489 17978
rect 15541 17926 24755 17978
rect 24807 17926 24819 17978
rect 24871 17926 24883 17978
rect 24935 17926 24947 17978
rect 24999 17926 25011 17978
rect 25063 17926 34277 17978
rect 34329 17926 34341 17978
rect 34393 17926 34405 17978
rect 34457 17926 34469 17978
rect 34521 17926 34533 17978
rect 34585 17926 39192 17978
rect 1104 17904 39192 17926
rect 22922 17864 22928 17876
rect 2746 17836 22928 17864
rect 1762 17688 1768 17740
rect 1820 17728 1826 17740
rect 2746 17728 2774 17836
rect 22922 17824 22928 17836
rect 22980 17824 22986 17876
rect 25774 17824 25780 17876
rect 25832 17864 25838 17876
rect 25961 17867 26019 17873
rect 25961 17864 25973 17867
rect 25832 17836 25973 17864
rect 25832 17824 25838 17836
rect 25961 17833 25973 17836
rect 26007 17833 26019 17867
rect 25961 17827 26019 17833
rect 26142 17824 26148 17876
rect 26200 17824 26206 17876
rect 27614 17864 27620 17876
rect 26252 17836 27620 17864
rect 21082 17756 21088 17808
rect 21140 17756 21146 17808
rect 24581 17799 24639 17805
rect 24581 17765 24593 17799
rect 24627 17765 24639 17799
rect 26252 17796 26280 17836
rect 27614 17824 27620 17836
rect 27672 17824 27678 17876
rect 28718 17824 28724 17876
rect 28776 17864 28782 17876
rect 29086 17864 29092 17876
rect 28776 17836 29092 17864
rect 28776 17824 28782 17836
rect 29086 17824 29092 17836
rect 29144 17824 29150 17876
rect 24581 17759 24639 17765
rect 24688 17768 26280 17796
rect 26697 17799 26755 17805
rect 1820 17700 2774 17728
rect 15933 17731 15991 17737
rect 1820 17688 1826 17700
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 18046 17728 18052 17740
rect 15979 17700 18052 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 18046 17688 18052 17700
rect 18104 17688 18110 17740
rect 21729 17731 21787 17737
rect 21729 17697 21741 17731
rect 21775 17728 21787 17731
rect 21775 17700 22232 17728
rect 21775 17697 21787 17700
rect 21729 17691 21787 17697
rect 2038 17620 2044 17672
rect 2096 17620 2102 17672
rect 2685 17663 2743 17669
rect 2685 17629 2697 17663
rect 2731 17660 2743 17663
rect 6638 17660 6644 17672
rect 2731 17632 6644 17660
rect 2731 17629 2743 17632
rect 2685 17623 2743 17629
rect 6638 17620 6644 17632
rect 6696 17620 6702 17672
rect 14090 17620 14096 17672
rect 14148 17660 14154 17672
rect 15654 17660 15660 17672
rect 14148 17632 15660 17660
rect 14148 17620 14154 17632
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 20257 17663 20315 17669
rect 20257 17629 20269 17663
rect 20303 17660 20315 17663
rect 20346 17660 20352 17672
rect 20303 17632 20352 17660
rect 20303 17629 20315 17632
rect 20257 17623 20315 17629
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20530 17620 20536 17672
rect 20588 17660 20594 17672
rect 22094 17662 22100 17672
rect 22066 17660 22100 17662
rect 20588 17632 22100 17660
rect 20588 17620 20594 17632
rect 22094 17620 22100 17632
rect 22152 17620 22158 17672
rect 22204 17660 22232 17700
rect 22278 17688 22284 17740
rect 22336 17688 22342 17740
rect 22557 17731 22615 17737
rect 22557 17697 22569 17731
rect 22603 17728 22615 17731
rect 24596 17728 24624 17759
rect 22603 17700 24624 17728
rect 22603 17697 22615 17700
rect 22557 17691 22615 17697
rect 22204 17632 22324 17660
rect 17310 17592 17316 17604
rect 17158 17564 17316 17592
rect 17310 17552 17316 17564
rect 17368 17552 17374 17604
rect 21082 17552 21088 17604
rect 21140 17592 21146 17604
rect 21545 17595 21603 17601
rect 21545 17592 21557 17595
rect 21140 17564 21557 17592
rect 21140 17552 21146 17564
rect 21545 17561 21557 17564
rect 21591 17561 21603 17595
rect 21545 17555 21603 17561
rect 2133 17527 2191 17533
rect 2133 17493 2145 17527
rect 2179 17524 2191 17527
rect 2406 17524 2412 17536
rect 2179 17496 2412 17524
rect 2179 17493 2191 17496
rect 2133 17487 2191 17493
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 2774 17484 2780 17536
rect 2832 17484 2838 17536
rect 17405 17527 17463 17533
rect 17405 17493 17417 17527
rect 17451 17524 17463 17527
rect 17494 17524 17500 17536
rect 17451 17496 17500 17524
rect 17451 17493 17463 17496
rect 17405 17487 17463 17493
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 19794 17484 19800 17536
rect 19852 17524 19858 17536
rect 19978 17524 19984 17536
rect 19852 17496 19984 17524
rect 19852 17484 19858 17496
rect 19978 17484 19984 17496
rect 20036 17524 20042 17536
rect 20349 17527 20407 17533
rect 20349 17524 20361 17527
rect 20036 17496 20361 17524
rect 20036 17484 20042 17496
rect 20349 17493 20361 17496
rect 20395 17493 20407 17527
rect 20349 17487 20407 17493
rect 21453 17527 21511 17533
rect 21453 17493 21465 17527
rect 21499 17524 21511 17527
rect 21726 17524 21732 17536
rect 21499 17496 21732 17524
rect 21499 17493 21511 17496
rect 21453 17487 21511 17493
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 22296 17524 22324 17632
rect 23658 17620 23664 17672
rect 23716 17620 23722 17672
rect 24688 17660 24716 17768
rect 26697 17765 26709 17799
rect 26743 17796 26755 17799
rect 27154 17796 27160 17808
rect 26743 17768 27160 17796
rect 26743 17765 26755 17768
rect 26697 17759 26755 17765
rect 27154 17756 27160 17768
rect 27212 17756 27218 17808
rect 28442 17756 28448 17808
rect 28500 17796 28506 17808
rect 30558 17796 30564 17808
rect 28500 17768 30564 17796
rect 28500 17756 28506 17768
rect 30558 17756 30564 17768
rect 30616 17756 30622 17808
rect 32490 17756 32496 17808
rect 32548 17796 32554 17808
rect 33962 17796 33968 17808
rect 32548 17768 33968 17796
rect 32548 17756 32554 17768
rect 33962 17756 33968 17768
rect 34020 17756 34026 17808
rect 25222 17688 25228 17740
rect 25280 17688 25286 17740
rect 27338 17688 27344 17740
rect 27396 17728 27402 17740
rect 31018 17728 31024 17740
rect 27396 17700 31024 17728
rect 27396 17688 27402 17700
rect 31018 17688 31024 17700
rect 31076 17688 31082 17740
rect 31294 17688 31300 17740
rect 31352 17688 31358 17740
rect 31754 17688 31760 17740
rect 31812 17728 31818 17740
rect 33045 17731 33103 17737
rect 33045 17728 33057 17731
rect 31812 17700 33057 17728
rect 31812 17688 31818 17700
rect 33045 17697 33057 17700
rect 33091 17697 33103 17731
rect 33045 17691 33103 17697
rect 34606 17688 34612 17740
rect 34664 17728 34670 17740
rect 35894 17728 35900 17740
rect 34664 17700 35900 17728
rect 34664 17688 34670 17700
rect 35894 17688 35900 17700
rect 35952 17688 35958 17740
rect 23860 17632 24716 17660
rect 23860 17524 23888 17632
rect 24946 17620 24952 17672
rect 25004 17620 25010 17672
rect 27157 17663 27215 17669
rect 27157 17629 27169 17663
rect 27203 17660 27215 17663
rect 27246 17660 27252 17672
rect 27203 17632 27252 17660
rect 27203 17629 27215 17632
rect 27157 17623 27215 17629
rect 27246 17620 27252 17632
rect 27304 17620 27310 17672
rect 29733 17663 29791 17669
rect 29733 17629 29745 17663
rect 29779 17660 29791 17663
rect 30190 17660 30196 17672
rect 29779 17632 30196 17660
rect 29779 17629 29791 17632
rect 29733 17623 29791 17629
rect 30190 17620 30196 17632
rect 30248 17620 30254 17672
rect 30558 17620 30564 17672
rect 30616 17660 30622 17672
rect 30616 17632 31064 17660
rect 30616 17620 30622 17632
rect 25041 17595 25099 17601
rect 25041 17592 25053 17595
rect 24044 17564 25053 17592
rect 24044 17533 24072 17564
rect 25041 17561 25053 17564
rect 25087 17592 25099 17595
rect 25777 17595 25835 17601
rect 25777 17592 25789 17595
rect 25087 17564 25789 17592
rect 25087 17561 25099 17564
rect 25041 17555 25099 17561
rect 25777 17561 25789 17564
rect 25823 17561 25835 17595
rect 25777 17555 25835 17561
rect 25958 17552 25964 17604
rect 26016 17601 26022 17604
rect 26016 17595 26035 17601
rect 26023 17561 26035 17595
rect 26016 17555 26035 17561
rect 26697 17595 26755 17601
rect 26697 17561 26709 17595
rect 26743 17592 26755 17595
rect 26878 17592 26884 17604
rect 26743 17564 26884 17592
rect 26743 17561 26755 17564
rect 26697 17555 26755 17561
rect 26016 17552 26022 17555
rect 26878 17552 26884 17564
rect 26936 17552 26942 17604
rect 30650 17592 30656 17604
rect 27264 17564 30656 17592
rect 27264 17533 27292 17564
rect 30650 17552 30656 17564
rect 30708 17552 30714 17604
rect 31036 17592 31064 17632
rect 32766 17620 32772 17672
rect 32824 17660 32830 17672
rect 32824 17632 33088 17660
rect 32824 17620 32830 17632
rect 33060 17592 33088 17632
rect 33134 17620 33140 17672
rect 33192 17660 33198 17672
rect 33781 17663 33839 17669
rect 33781 17660 33793 17663
rect 33192 17632 33793 17660
rect 33192 17620 33198 17632
rect 33781 17629 33793 17632
rect 33827 17660 33839 17663
rect 37182 17660 37188 17672
rect 33827 17632 37188 17660
rect 33827 17629 33839 17632
rect 33781 17623 33839 17629
rect 37182 17620 37188 17632
rect 37240 17620 37246 17672
rect 35158 17592 35164 17604
rect 31036 17564 31340 17592
rect 32522 17564 32812 17592
rect 33060 17564 35164 17592
rect 22296 17496 23888 17524
rect 24029 17527 24087 17533
rect 24029 17493 24041 17527
rect 24075 17493 24087 17527
rect 24029 17487 24087 17493
rect 27249 17527 27307 17533
rect 27249 17493 27261 17527
rect 27295 17493 27307 17527
rect 27249 17487 27307 17493
rect 27430 17484 27436 17536
rect 27488 17484 27494 17536
rect 27522 17484 27528 17536
rect 27580 17524 27586 17536
rect 29825 17527 29883 17533
rect 29825 17524 29837 17527
rect 27580 17496 29837 17524
rect 27580 17484 27586 17496
rect 29825 17493 29837 17496
rect 29871 17493 29883 17527
rect 29825 17487 29883 17493
rect 30282 17484 30288 17536
rect 30340 17524 30346 17536
rect 31202 17524 31208 17536
rect 30340 17496 31208 17524
rect 30340 17484 30346 17496
rect 31202 17484 31208 17496
rect 31260 17484 31266 17536
rect 31312 17524 31340 17564
rect 32582 17524 32588 17536
rect 31312 17496 32588 17524
rect 32582 17484 32588 17496
rect 32640 17484 32646 17536
rect 32784 17524 32812 17564
rect 35158 17552 35164 17564
rect 35216 17552 35222 17604
rect 33873 17527 33931 17533
rect 33873 17524 33885 17527
rect 32784 17496 33885 17524
rect 33873 17493 33885 17496
rect 33919 17493 33931 17527
rect 33873 17487 33931 17493
rect 1104 17434 39352 17456
rect 1104 17382 10472 17434
rect 10524 17382 10536 17434
rect 10588 17382 10600 17434
rect 10652 17382 10664 17434
rect 10716 17382 10728 17434
rect 10780 17382 19994 17434
rect 20046 17382 20058 17434
rect 20110 17382 20122 17434
rect 20174 17382 20186 17434
rect 20238 17382 20250 17434
rect 20302 17382 29516 17434
rect 29568 17382 29580 17434
rect 29632 17382 29644 17434
rect 29696 17382 29708 17434
rect 29760 17382 29772 17434
rect 29824 17382 39038 17434
rect 39090 17382 39102 17434
rect 39154 17382 39166 17434
rect 39218 17382 39230 17434
rect 39282 17382 39294 17434
rect 39346 17382 39352 17434
rect 1104 17360 39352 17382
rect 6822 17280 6828 17332
rect 6880 17320 6886 17332
rect 7374 17320 7380 17332
rect 6880 17292 7380 17320
rect 6880 17280 6886 17292
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 7653 17323 7711 17329
rect 7653 17289 7665 17323
rect 7699 17320 7711 17323
rect 7699 17292 12434 17320
rect 7699 17289 7711 17292
rect 7653 17283 7711 17289
rect 5261 17255 5319 17261
rect 5261 17221 5273 17255
rect 5307 17252 5319 17255
rect 7742 17252 7748 17264
rect 5307 17224 7748 17252
rect 5307 17221 5319 17224
rect 5261 17215 5319 17221
rect 7742 17212 7748 17224
rect 7800 17252 7806 17264
rect 9490 17252 9496 17264
rect 7800 17224 9496 17252
rect 7800 17212 7806 17224
rect 9490 17212 9496 17224
rect 9548 17212 9554 17264
rect 12406 17252 12434 17292
rect 13630 17280 13636 17332
rect 13688 17320 13694 17332
rect 13688 17292 14504 17320
rect 13688 17280 13694 17292
rect 14369 17255 14427 17261
rect 14369 17252 14381 17255
rect 12406 17224 14381 17252
rect 14369 17221 14381 17224
rect 14415 17221 14427 17255
rect 14476 17252 14504 17292
rect 19794 17280 19800 17332
rect 19852 17320 19858 17332
rect 19852 17292 22094 17320
rect 19852 17280 19858 17292
rect 14476 17224 14858 17252
rect 14369 17215 14427 17221
rect 17126 17212 17132 17264
rect 17184 17212 17190 17264
rect 18138 17212 18144 17264
rect 18196 17212 18202 17264
rect 22066 17252 22094 17292
rect 23934 17280 23940 17332
rect 23992 17280 23998 17332
rect 24118 17280 24124 17332
rect 24176 17320 24182 17332
rect 24176 17292 25912 17320
rect 24176 17280 24182 17292
rect 23201 17255 23259 17261
rect 22066 17224 23152 17252
rect 1578 17144 1584 17196
rect 1636 17144 1642 17196
rect 3970 17144 3976 17196
rect 4028 17144 4034 17196
rect 5166 17144 5172 17196
rect 5224 17144 5230 17196
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8076 17156 12434 17184
rect 8076 17144 8082 17156
rect 2222 17076 2228 17128
rect 2280 17116 2286 17128
rect 2593 17119 2651 17125
rect 2593 17116 2605 17119
rect 2280 17088 2605 17116
rect 2280 17076 2286 17088
rect 2593 17085 2605 17088
rect 2639 17085 2651 17119
rect 2593 17079 2651 17085
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 4338 17116 4344 17128
rect 2915 17088 4344 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 4338 17076 4344 17088
rect 4396 17076 4402 17128
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17085 5411 17119
rect 5353 17079 5411 17085
rect 5074 17008 5080 17060
rect 5132 17048 5138 17060
rect 5368 17048 5396 17079
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 5592 17088 8125 17116
rect 5592 17076 5598 17088
rect 8113 17085 8125 17088
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 10870 17116 10876 17128
rect 8251 17088 10876 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 10870 17076 10876 17088
rect 10928 17116 10934 17128
rect 11882 17116 11888 17128
rect 10928 17088 11888 17116
rect 10928 17076 10934 17088
rect 11882 17076 11888 17088
rect 11940 17076 11946 17128
rect 12406 17116 12434 17156
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 14090 17184 14096 17196
rect 13228 17156 14096 17184
rect 13228 17144 13234 17156
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 15654 17144 15660 17196
rect 15712 17184 15718 17196
rect 16850 17184 16856 17196
rect 15712 17156 16856 17184
rect 15712 17144 15718 17156
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 22557 17187 22615 17193
rect 16117 17119 16175 17125
rect 12406 17088 14228 17116
rect 5132 17020 5396 17048
rect 5132 17008 5138 17020
rect 1673 16983 1731 16989
rect 1673 16949 1685 16983
rect 1719 16980 1731 16983
rect 1854 16980 1860 16992
rect 1719 16952 1860 16980
rect 1719 16949 1731 16952
rect 1673 16943 1731 16949
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 4341 16983 4399 16989
rect 4341 16949 4353 16983
rect 4387 16980 4399 16983
rect 4430 16980 4436 16992
rect 4387 16952 4436 16980
rect 4387 16949 4399 16952
rect 4341 16943 4399 16949
rect 4430 16940 4436 16952
rect 4488 16940 4494 16992
rect 4798 16940 4804 16992
rect 4856 16940 4862 16992
rect 5350 16940 5356 16992
rect 5408 16980 5414 16992
rect 6822 16980 6828 16992
rect 5408 16952 6828 16980
rect 5408 16940 5414 16952
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 14200 16980 14228 17088
rect 16117 17085 16129 17119
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 16132 16980 16160 17079
rect 16482 17076 16488 17128
rect 16540 17116 16546 17128
rect 18782 17116 18788 17128
rect 16540 17088 18788 17116
rect 16540 17076 16546 17088
rect 18782 17076 18788 17088
rect 18840 17116 18846 17128
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 18840 17088 18889 17116
rect 18840 17076 18846 17088
rect 18877 17085 18889 17088
rect 18923 17085 18935 17119
rect 18877 17079 18935 17085
rect 19337 17119 19395 17125
rect 19337 17085 19349 17119
rect 19383 17085 19395 17119
rect 19337 17079 19395 17085
rect 19613 17119 19671 17125
rect 19613 17085 19625 17119
rect 19659 17116 19671 17119
rect 20732 17116 20760 17170
rect 22557 17153 22569 17187
rect 22603 17184 22615 17187
rect 22830 17184 22836 17196
rect 22603 17156 22836 17184
rect 22603 17153 22615 17156
rect 22557 17147 22615 17153
rect 22830 17144 22836 17156
rect 22888 17144 22894 17196
rect 20806 17116 20812 17128
rect 19659 17088 20668 17116
rect 20732 17088 20812 17116
rect 19659 17085 19671 17088
rect 19613 17079 19671 17085
rect 14200 16952 16160 16980
rect 19352 16980 19380 17079
rect 20640 17048 20668 17088
rect 20806 17076 20812 17088
rect 20864 17076 20870 17128
rect 23124 17116 23152 17224
rect 23201 17221 23213 17255
rect 23247 17252 23259 17255
rect 23382 17252 23388 17264
rect 23247 17224 23388 17252
rect 23247 17221 23259 17224
rect 23201 17215 23259 17221
rect 23382 17212 23388 17224
rect 23440 17212 23446 17264
rect 24578 17212 24584 17264
rect 24636 17252 24642 17264
rect 25225 17255 25283 17261
rect 25225 17252 25237 17255
rect 24636 17224 25237 17252
rect 24636 17212 24642 17224
rect 25225 17221 25237 17224
rect 25271 17221 25283 17255
rect 25225 17215 25283 17221
rect 23400 17184 23428 17212
rect 23842 17184 23848 17196
rect 23400 17156 23848 17184
rect 23842 17144 23848 17156
rect 23900 17144 23906 17196
rect 24486 17144 24492 17196
rect 24544 17144 24550 17196
rect 25884 17193 25912 17292
rect 26326 17280 26332 17332
rect 26384 17320 26390 17332
rect 26421 17323 26479 17329
rect 26421 17320 26433 17323
rect 26384 17292 26433 17320
rect 26384 17280 26390 17292
rect 26421 17289 26433 17292
rect 26467 17289 26479 17323
rect 26421 17283 26479 17289
rect 30101 17323 30159 17329
rect 30101 17289 30113 17323
rect 30147 17320 30159 17323
rect 32766 17320 32772 17332
rect 30147 17292 32772 17320
rect 30147 17289 30159 17292
rect 30101 17283 30159 17289
rect 32766 17280 32772 17292
rect 32824 17280 32830 17332
rect 32950 17280 32956 17332
rect 33008 17280 33014 17332
rect 38562 17320 38568 17332
rect 33060 17292 38568 17320
rect 25976 17224 26280 17252
rect 25869 17187 25927 17193
rect 25869 17153 25881 17187
rect 25915 17153 25927 17187
rect 25869 17147 25927 17153
rect 25976 17116 26004 17224
rect 26050 17144 26056 17196
rect 26108 17144 26114 17196
rect 26252 17193 26280 17224
rect 26694 17212 26700 17264
rect 26752 17252 26758 17264
rect 27249 17255 27307 17261
rect 27249 17252 27261 17255
rect 26752 17224 27261 17252
rect 26752 17212 26758 17224
rect 27249 17221 27261 17224
rect 27295 17221 27307 17255
rect 27249 17215 27307 17221
rect 27430 17212 27436 17264
rect 27488 17252 27494 17264
rect 27488 17224 30972 17252
rect 27488 17212 27494 17224
rect 26145 17187 26203 17193
rect 26145 17153 26157 17187
rect 26191 17153 26203 17187
rect 26145 17147 26203 17153
rect 26237 17187 26295 17193
rect 26237 17153 26249 17187
rect 26283 17184 26295 17187
rect 28350 17184 28356 17196
rect 26283 17156 28356 17184
rect 26283 17153 26295 17156
rect 26237 17147 26295 17153
rect 23124 17088 26004 17116
rect 26160 17116 26188 17147
rect 28350 17144 28356 17156
rect 28408 17144 28414 17196
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 30009 17187 30067 17193
rect 30009 17184 30021 17187
rect 29052 17156 30021 17184
rect 29052 17144 29058 17156
rect 30009 17153 30021 17156
rect 30055 17184 30067 17187
rect 30098 17184 30104 17196
rect 30055 17156 30104 17184
rect 30055 17153 30067 17156
rect 30009 17147 30067 17153
rect 30098 17144 30104 17156
rect 30156 17144 30162 17196
rect 30374 17144 30380 17196
rect 30432 17184 30438 17196
rect 30558 17184 30564 17196
rect 30432 17156 30564 17184
rect 30432 17144 30438 17156
rect 30558 17144 30564 17156
rect 30616 17144 30622 17196
rect 30834 17144 30840 17196
rect 30892 17144 30898 17196
rect 30944 17184 30972 17224
rect 31018 17212 31024 17264
rect 31076 17252 31082 17264
rect 31573 17255 31631 17261
rect 31573 17252 31585 17255
rect 31076 17224 31585 17252
rect 31076 17212 31082 17224
rect 31573 17221 31585 17224
rect 31619 17221 31631 17255
rect 31573 17215 31631 17221
rect 32582 17212 32588 17264
rect 32640 17212 32646 17264
rect 32677 17255 32735 17261
rect 32677 17221 32689 17255
rect 32723 17252 32735 17255
rect 33060 17252 33088 17292
rect 38562 17280 38568 17292
rect 38620 17280 38626 17332
rect 32723 17224 33088 17252
rect 32723 17221 32735 17224
rect 32677 17215 32735 17221
rect 33962 17212 33968 17264
rect 34020 17252 34026 17264
rect 34241 17255 34299 17261
rect 34241 17252 34253 17255
rect 34020 17224 34253 17252
rect 34020 17212 34026 17224
rect 34241 17221 34253 17224
rect 34287 17221 34299 17255
rect 34241 17215 34299 17221
rect 34330 17212 34336 17264
rect 34388 17252 34394 17264
rect 35437 17255 35495 17261
rect 35437 17252 35449 17255
rect 34388 17224 35449 17252
rect 34388 17212 34394 17224
rect 35437 17221 35449 17224
rect 35483 17252 35495 17255
rect 35710 17252 35716 17264
rect 35483 17224 35716 17252
rect 35483 17221 35495 17224
rect 35437 17215 35495 17221
rect 35710 17212 35716 17224
rect 35768 17212 35774 17264
rect 32309 17187 32367 17193
rect 32309 17184 32321 17187
rect 30944 17156 32321 17184
rect 32309 17153 32321 17156
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 32402 17187 32460 17193
rect 32402 17153 32414 17187
rect 32448 17153 32460 17187
rect 32815 17187 32873 17193
rect 32815 17184 32827 17187
rect 32402 17147 32460 17153
rect 32600 17156 32827 17184
rect 29178 17116 29184 17128
rect 26160 17088 29184 17116
rect 29178 17076 29184 17088
rect 29236 17116 29242 17128
rect 29730 17116 29736 17128
rect 29236 17088 29736 17116
rect 29236 17076 29242 17088
rect 29730 17076 29736 17088
rect 29788 17076 29794 17128
rect 29914 17076 29920 17128
rect 29972 17116 29978 17128
rect 30285 17119 30343 17125
rect 30285 17116 30297 17119
rect 29972 17088 30297 17116
rect 29972 17076 29978 17088
rect 30285 17085 30297 17088
rect 30331 17116 30343 17119
rect 31570 17116 31576 17128
rect 30331 17088 31576 17116
rect 30331 17085 30343 17088
rect 30285 17079 30343 17085
rect 31570 17076 31576 17088
rect 31628 17076 31634 17128
rect 31662 17076 31668 17128
rect 31720 17116 31726 17128
rect 32416 17116 32444 17147
rect 31720 17088 32444 17116
rect 31720 17076 31726 17088
rect 21634 17048 21640 17060
rect 20640 17020 21640 17048
rect 21634 17008 21640 17020
rect 21692 17008 21698 17060
rect 29362 17008 29368 17060
rect 29420 17048 29426 17060
rect 29420 17020 30236 17048
rect 29420 17008 29426 17020
rect 20990 16980 20996 16992
rect 19352 16952 20996 16980
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 21085 16983 21143 16989
rect 21085 16949 21097 16983
rect 21131 16980 21143 16983
rect 21542 16980 21548 16992
rect 21131 16952 21548 16980
rect 21131 16949 21143 16952
rect 21085 16943 21143 16949
rect 21542 16940 21548 16952
rect 21600 16940 21606 16992
rect 27154 16940 27160 16992
rect 27212 16980 27218 16992
rect 27341 16983 27399 16989
rect 27341 16980 27353 16983
rect 27212 16952 27353 16980
rect 27212 16940 27218 16952
rect 27341 16949 27353 16952
rect 27387 16949 27399 16983
rect 27341 16943 27399 16949
rect 27614 16940 27620 16992
rect 27672 16980 27678 16992
rect 27982 16980 27988 16992
rect 27672 16952 27988 16980
rect 27672 16940 27678 16952
rect 27982 16940 27988 16952
rect 28040 16940 28046 16992
rect 29641 16983 29699 16989
rect 29641 16949 29653 16983
rect 29687 16980 29699 16983
rect 30098 16980 30104 16992
rect 29687 16952 30104 16980
rect 29687 16949 29699 16952
rect 29641 16943 29699 16949
rect 30098 16940 30104 16952
rect 30156 16940 30162 16992
rect 30208 16980 30236 17020
rect 30374 17008 30380 17060
rect 30432 17048 30438 17060
rect 32600 17048 32628 17156
rect 32815 17153 32827 17156
rect 32861 17184 32873 17187
rect 32861 17156 34008 17184
rect 32861 17153 32873 17156
rect 32815 17147 32873 17153
rect 32674 17076 32680 17128
rect 32732 17116 32738 17128
rect 33980 17116 34008 17156
rect 34146 17144 34152 17196
rect 34204 17144 34210 17196
rect 34256 17156 34468 17184
rect 34256 17116 34284 17156
rect 32732 17088 33916 17116
rect 33980 17088 34284 17116
rect 32732 17076 32738 17088
rect 33781 17051 33839 17057
rect 33781 17048 33793 17051
rect 30432 17020 32628 17048
rect 32876 17020 33793 17048
rect 30432 17008 30438 17020
rect 32876 16980 32904 17020
rect 33781 17017 33793 17020
rect 33827 17017 33839 17051
rect 33888 17048 33916 17088
rect 34330 17076 34336 17128
rect 34388 17076 34394 17128
rect 34440 17116 34468 17156
rect 34882 17144 34888 17196
rect 34940 17184 34946 17196
rect 35069 17187 35127 17193
rect 35069 17184 35081 17187
rect 34940 17156 35081 17184
rect 34940 17144 34946 17156
rect 35069 17153 35081 17156
rect 35115 17153 35127 17187
rect 35069 17147 35127 17153
rect 37366 17144 37372 17196
rect 37424 17184 37430 17196
rect 38473 17187 38531 17193
rect 38473 17184 38485 17187
rect 37424 17156 38485 17184
rect 37424 17144 37430 17156
rect 38473 17153 38485 17156
rect 38519 17153 38531 17187
rect 38473 17147 38531 17153
rect 35250 17116 35256 17128
rect 34440 17088 35256 17116
rect 35250 17076 35256 17088
rect 35308 17076 35314 17128
rect 36446 17048 36452 17060
rect 33888 17020 36452 17048
rect 33781 17011 33839 17017
rect 36446 17008 36452 17020
rect 36504 17008 36510 17060
rect 38654 17008 38660 17060
rect 38712 17008 38718 17060
rect 30208 16952 32904 16980
rect 1104 16890 39192 16912
rect 1104 16838 5711 16890
rect 5763 16838 5775 16890
rect 5827 16838 5839 16890
rect 5891 16838 5903 16890
rect 5955 16838 5967 16890
rect 6019 16838 15233 16890
rect 15285 16838 15297 16890
rect 15349 16838 15361 16890
rect 15413 16838 15425 16890
rect 15477 16838 15489 16890
rect 15541 16838 24755 16890
rect 24807 16838 24819 16890
rect 24871 16838 24883 16890
rect 24935 16838 24947 16890
rect 24999 16838 25011 16890
rect 25063 16838 34277 16890
rect 34329 16838 34341 16890
rect 34393 16838 34405 16890
rect 34457 16838 34469 16890
rect 34521 16838 34533 16890
rect 34585 16838 39192 16890
rect 1104 16816 39192 16838
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16776 2007 16779
rect 5350 16776 5356 16788
rect 1995 16748 5356 16776
rect 1995 16745 2007 16748
rect 1949 16739 2007 16745
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 5442 16736 5448 16788
rect 5500 16776 5506 16788
rect 5994 16776 6000 16788
rect 5500 16748 6000 16776
rect 5500 16736 5506 16748
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 12526 16736 12532 16788
rect 12584 16776 12590 16788
rect 12805 16779 12863 16785
rect 12805 16776 12817 16779
rect 12584 16748 12817 16776
rect 12584 16736 12590 16748
rect 12805 16745 12817 16748
rect 12851 16745 12863 16779
rect 12805 16739 12863 16745
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 17218 16776 17224 16788
rect 13872 16748 17224 16776
rect 13872 16736 13878 16748
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 17954 16736 17960 16788
rect 18012 16776 18018 16788
rect 18138 16776 18144 16788
rect 18012 16748 18144 16776
rect 18012 16736 18018 16748
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 20990 16736 20996 16788
rect 21048 16776 21054 16788
rect 22278 16776 22284 16788
rect 21048 16748 22284 16776
rect 21048 16736 21054 16748
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 26602 16736 26608 16788
rect 26660 16736 26666 16788
rect 34348 16748 35204 16776
rect 12989 16711 13047 16717
rect 12989 16677 13001 16711
rect 13035 16708 13047 16711
rect 15378 16708 15384 16720
rect 13035 16680 15384 16708
rect 13035 16677 13047 16680
rect 12989 16671 13047 16677
rect 15378 16668 15384 16680
rect 15436 16668 15442 16720
rect 25130 16708 25136 16720
rect 23768 16680 25136 16708
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 4801 16643 4859 16649
rect 4801 16640 4813 16643
rect 4672 16612 4813 16640
rect 4672 16600 4678 16612
rect 4801 16609 4813 16612
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 4890 16600 4896 16652
rect 4948 16600 4954 16652
rect 11790 16600 11796 16652
rect 11848 16640 11854 16652
rect 12250 16640 12256 16652
rect 11848 16612 12256 16640
rect 11848 16600 11854 16612
rect 12250 16600 12256 16612
rect 12308 16640 12314 16652
rect 13814 16640 13820 16652
rect 12308 16612 13820 16640
rect 12308 16600 12314 16612
rect 2038 16532 2044 16584
rect 2096 16572 2102 16584
rect 2593 16575 2651 16581
rect 2593 16572 2605 16575
rect 2096 16544 2605 16572
rect 2096 16532 2102 16544
rect 2593 16541 2605 16544
rect 2639 16572 2651 16575
rect 3142 16572 3148 16584
rect 2639 16544 3148 16572
rect 2639 16541 2651 16544
rect 2593 16535 2651 16541
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 3237 16575 3295 16581
rect 3237 16541 3249 16575
rect 3283 16572 3295 16575
rect 5537 16575 5595 16581
rect 5537 16572 5549 16575
rect 3283 16544 5549 16572
rect 3283 16541 3295 16544
rect 3237 16535 3295 16541
rect 5537 16541 5549 16544
rect 5583 16572 5595 16575
rect 5626 16572 5632 16584
rect 5583 16544 5632 16572
rect 5583 16541 5595 16544
rect 5537 16535 5595 16541
rect 5626 16532 5632 16544
rect 5684 16572 5690 16584
rect 6181 16575 6239 16581
rect 6181 16572 6193 16575
rect 5684 16544 6193 16572
rect 5684 16532 5690 16544
rect 6181 16541 6193 16544
rect 6227 16541 6239 16575
rect 6181 16535 6239 16541
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 9306 16572 9312 16584
rect 7800 16544 9312 16572
rect 7800 16532 7806 16544
rect 9306 16532 9312 16544
rect 9364 16572 9370 16584
rect 13556 16581 13584 16612
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 15930 16640 15936 16652
rect 14660 16612 15936 16640
rect 13541 16575 13599 16581
rect 9364 16547 12864 16572
rect 9364 16544 12909 16547
rect 9364 16532 9370 16544
rect 12836 16541 12909 16544
rect 934 16464 940 16516
rect 992 16504 998 16516
rect 1673 16507 1731 16513
rect 1673 16504 1685 16507
rect 992 16476 1685 16504
rect 992 16464 998 16476
rect 1673 16473 1685 16476
rect 1719 16473 1731 16507
rect 1673 16467 1731 16473
rect 12250 16464 12256 16516
rect 12308 16504 12314 16516
rect 12621 16507 12679 16513
rect 12621 16504 12633 16507
rect 12308 16476 12633 16504
rect 12308 16464 12314 16476
rect 12621 16473 12633 16476
rect 12667 16473 12679 16507
rect 12836 16507 12863 16541
rect 12897 16516 12909 16541
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 13630 16532 13636 16584
rect 13688 16532 13694 16584
rect 14660 16581 14688 16612
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 17236 16612 17908 16640
rect 17236 16584 17264 16612
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16541 14703 16575
rect 14921 16575 14979 16581
rect 14921 16572 14933 16575
rect 14645 16535 14703 16541
rect 14752 16544 14933 16572
rect 12897 16507 12900 16516
rect 12836 16476 12900 16507
rect 12621 16467 12679 16473
rect 12894 16464 12900 16476
rect 12952 16464 12958 16516
rect 14550 16464 14556 16516
rect 14608 16504 14614 16516
rect 14752 16504 14780 16544
rect 14921 16541 14933 16544
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15013 16575 15071 16581
rect 15013 16541 15025 16575
rect 15059 16572 15071 16575
rect 15102 16572 15108 16584
rect 15059 16544 15108 16572
rect 15059 16541 15071 16544
rect 15013 16535 15071 16541
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 14608 16476 14780 16504
rect 14829 16507 14887 16513
rect 14608 16464 14614 16476
rect 14829 16473 14841 16507
rect 14875 16504 14887 16507
rect 15654 16504 15660 16516
rect 14875 16476 15660 16504
rect 14875 16473 14887 16476
rect 14829 16467 14887 16473
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 15764 16504 15792 16535
rect 17218 16532 17224 16584
rect 17276 16532 17282 16584
rect 17310 16532 17316 16584
rect 17368 16532 17374 16584
rect 17880 16581 17908 16612
rect 20990 16600 20996 16652
rect 21048 16600 21054 16652
rect 21269 16643 21327 16649
rect 21269 16609 21281 16643
rect 21315 16640 21327 16643
rect 23014 16640 23020 16652
rect 21315 16612 23020 16640
rect 21315 16609 21327 16612
rect 21269 16603 21327 16609
rect 23014 16600 23020 16612
rect 23072 16600 23078 16652
rect 23566 16600 23572 16652
rect 23624 16640 23630 16652
rect 23768 16649 23796 16680
rect 25130 16668 25136 16680
rect 25188 16708 25194 16720
rect 25188 16680 25820 16708
rect 25188 16668 25194 16680
rect 25792 16652 25820 16680
rect 30392 16680 30788 16708
rect 23661 16643 23719 16649
rect 23661 16640 23673 16643
rect 23624 16612 23673 16640
rect 23624 16600 23630 16612
rect 23661 16609 23673 16612
rect 23707 16609 23719 16643
rect 23661 16603 23719 16609
rect 23753 16643 23811 16649
rect 23753 16609 23765 16643
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 25314 16600 25320 16652
rect 25372 16600 25378 16652
rect 25774 16600 25780 16652
rect 25832 16640 25838 16652
rect 30392 16640 30420 16680
rect 25832 16612 30420 16640
rect 25832 16600 25838 16612
rect 30650 16600 30656 16652
rect 30708 16600 30714 16652
rect 30760 16649 30788 16680
rect 32858 16668 32864 16720
rect 32916 16708 32922 16720
rect 33045 16711 33103 16717
rect 33045 16708 33057 16711
rect 32916 16680 33057 16708
rect 32916 16668 32922 16680
rect 33045 16677 33057 16680
rect 33091 16677 33103 16711
rect 33045 16671 33103 16677
rect 33137 16711 33195 16717
rect 33137 16677 33149 16711
rect 33183 16708 33195 16711
rect 34348 16708 34376 16748
rect 33183 16680 34376 16708
rect 35176 16708 35204 16748
rect 35437 16711 35495 16717
rect 35437 16708 35449 16711
rect 35176 16680 35449 16708
rect 33183 16677 33195 16680
rect 33137 16671 33195 16677
rect 35437 16677 35449 16680
rect 35483 16677 35495 16711
rect 35437 16671 35495 16677
rect 30745 16643 30803 16649
rect 30745 16609 30757 16643
rect 30791 16640 30803 16643
rect 32674 16640 32680 16652
rect 30791 16612 32680 16640
rect 30791 16609 30803 16612
rect 30745 16603 30803 16609
rect 32674 16600 32680 16612
rect 32732 16600 32738 16652
rect 32769 16643 32827 16649
rect 32769 16609 32781 16643
rect 32815 16640 32827 16643
rect 35066 16640 35072 16652
rect 32815 16612 35072 16640
rect 32815 16609 32827 16612
rect 32769 16603 32827 16609
rect 35066 16600 35072 16612
rect 35124 16600 35130 16652
rect 35176 16612 35388 16640
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 23842 16532 23848 16584
rect 23900 16572 23906 16584
rect 26326 16572 26332 16584
rect 23900 16544 26332 16572
rect 23900 16532 23906 16544
rect 26326 16532 26332 16544
rect 26384 16572 26390 16584
rect 26605 16575 26663 16581
rect 26605 16572 26617 16575
rect 26384 16544 26617 16572
rect 26384 16532 26390 16544
rect 26605 16541 26617 16544
rect 26651 16541 26663 16575
rect 26605 16535 26663 16541
rect 27338 16532 27344 16584
rect 27396 16532 27402 16584
rect 28902 16532 28908 16584
rect 28960 16572 28966 16584
rect 30834 16572 30840 16584
rect 28960 16544 30840 16572
rect 28960 16532 28966 16544
rect 30834 16532 30840 16544
rect 30892 16572 30898 16584
rect 31389 16575 31447 16581
rect 31389 16572 31401 16575
rect 30892 16544 31401 16572
rect 30892 16532 30898 16544
rect 31389 16541 31401 16544
rect 31435 16541 31447 16575
rect 31389 16535 31447 16541
rect 31726 16544 33088 16572
rect 15764 16476 16160 16504
rect 2682 16396 2688 16448
rect 2740 16396 2746 16448
rect 3234 16396 3240 16448
rect 3292 16436 3298 16448
rect 3329 16439 3387 16445
rect 3329 16436 3341 16439
rect 3292 16408 3341 16436
rect 3292 16396 3298 16408
rect 3329 16405 3341 16408
rect 3375 16405 3387 16439
rect 3329 16399 3387 16405
rect 4338 16396 4344 16448
rect 4396 16396 4402 16448
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 4709 16439 4767 16445
rect 4709 16436 4721 16439
rect 4488 16408 4721 16436
rect 4488 16396 4494 16408
rect 4709 16405 4721 16408
rect 4755 16436 4767 16439
rect 4982 16436 4988 16448
rect 4755 16408 4988 16436
rect 4755 16405 4767 16408
rect 4709 16399 4767 16405
rect 4982 16396 4988 16408
rect 5040 16396 5046 16448
rect 5442 16396 5448 16448
rect 5500 16436 5506 16448
rect 5629 16439 5687 16445
rect 5629 16436 5641 16439
rect 5500 16408 5641 16436
rect 5500 16396 5506 16408
rect 5629 16405 5641 16408
rect 5675 16405 5687 16439
rect 5629 16399 5687 16405
rect 6273 16439 6331 16445
rect 6273 16405 6285 16439
rect 6319 16436 6331 16439
rect 12710 16436 12716 16448
rect 6319 16408 12716 16436
rect 6319 16405 6331 16408
rect 6273 16399 6331 16405
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 15197 16439 15255 16445
rect 15197 16405 15209 16439
rect 15243 16436 15255 16439
rect 16022 16436 16028 16448
rect 15243 16408 16028 16436
rect 15243 16405 15255 16408
rect 15197 16399 15255 16405
rect 16022 16396 16028 16408
rect 16080 16396 16086 16448
rect 16132 16436 16160 16476
rect 16298 16464 16304 16516
rect 16356 16464 16362 16516
rect 20714 16504 20720 16516
rect 16776 16476 20720 16504
rect 16776 16448 16804 16476
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 22278 16464 22284 16516
rect 22336 16464 22342 16516
rect 24486 16464 24492 16516
rect 24544 16504 24550 16516
rect 24581 16507 24639 16513
rect 24581 16504 24593 16507
rect 24544 16476 24593 16504
rect 24544 16464 24550 16476
rect 24581 16473 24593 16476
rect 24627 16473 24639 16507
rect 24581 16467 24639 16473
rect 16758 16436 16764 16448
rect 16132 16408 16764 16436
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 17954 16396 17960 16448
rect 18012 16396 18018 16448
rect 22738 16396 22744 16448
rect 22796 16396 22802 16448
rect 23198 16396 23204 16448
rect 23256 16396 23262 16448
rect 23569 16439 23627 16445
rect 23569 16405 23581 16439
rect 23615 16436 23627 16439
rect 23750 16436 23756 16448
rect 23615 16408 23756 16436
rect 23615 16405 23627 16408
rect 23569 16399 23627 16405
rect 23750 16396 23756 16408
rect 23808 16396 23814 16448
rect 24596 16436 24624 16467
rect 27614 16464 27620 16516
rect 27672 16464 27678 16516
rect 31726 16504 31754 16544
rect 28842 16476 31754 16504
rect 32217 16507 32275 16513
rect 32217 16473 32229 16507
rect 32263 16504 32275 16507
rect 32306 16504 32312 16516
rect 32263 16476 32312 16504
rect 32263 16473 32275 16476
rect 32217 16467 32275 16473
rect 32306 16464 32312 16476
rect 32364 16504 32370 16516
rect 32950 16504 32956 16516
rect 32364 16476 32956 16504
rect 32364 16464 32370 16476
rect 32950 16464 32956 16476
rect 33008 16464 33014 16516
rect 33060 16504 33088 16544
rect 33226 16532 33232 16584
rect 33284 16532 33290 16584
rect 33502 16532 33508 16584
rect 33560 16532 33566 16584
rect 33962 16532 33968 16584
rect 34020 16572 34026 16584
rect 34149 16575 34207 16581
rect 34149 16572 34161 16575
rect 34020 16544 34161 16572
rect 34020 16532 34026 16544
rect 34149 16541 34161 16544
rect 34195 16541 34207 16575
rect 34149 16535 34207 16541
rect 34885 16575 34943 16581
rect 34885 16541 34897 16575
rect 34931 16572 34943 16575
rect 35176 16572 35204 16612
rect 34931 16544 35204 16572
rect 34931 16541 34943 16544
rect 34885 16535 34943 16541
rect 35250 16532 35256 16584
rect 35308 16532 35314 16584
rect 35360 16572 35388 16612
rect 35526 16572 35532 16584
rect 35360 16544 35532 16572
rect 35526 16532 35532 16544
rect 35584 16532 35590 16584
rect 35897 16575 35955 16581
rect 35897 16541 35909 16575
rect 35943 16572 35955 16575
rect 36541 16575 36599 16581
rect 36541 16572 36553 16575
rect 35943 16544 36553 16572
rect 35943 16541 35955 16544
rect 35897 16535 35955 16541
rect 36541 16541 36553 16544
rect 36587 16572 36599 16575
rect 36630 16572 36636 16584
rect 36587 16544 36636 16572
rect 36587 16541 36599 16544
rect 36541 16535 36599 16541
rect 36630 16532 36636 16544
rect 36688 16532 36694 16584
rect 34241 16507 34299 16513
rect 34241 16504 34253 16507
rect 33060 16476 34253 16504
rect 34241 16473 34253 16476
rect 34287 16473 34299 16507
rect 34241 16467 34299 16473
rect 34330 16464 34336 16516
rect 34388 16504 34394 16516
rect 35069 16507 35127 16513
rect 35069 16504 35081 16507
rect 34388 16476 35081 16504
rect 34388 16464 34394 16476
rect 35069 16473 35081 16476
rect 35115 16473 35127 16507
rect 35069 16467 35127 16473
rect 35158 16464 35164 16516
rect 35216 16464 35222 16516
rect 25222 16436 25228 16448
rect 24596 16408 25228 16436
rect 25222 16396 25228 16408
rect 25280 16436 25286 16448
rect 28902 16436 28908 16448
rect 25280 16408 28908 16436
rect 25280 16396 25286 16408
rect 28902 16396 28908 16408
rect 28960 16396 28966 16448
rect 28994 16396 29000 16448
rect 29052 16436 29058 16448
rect 29089 16439 29147 16445
rect 29089 16436 29101 16439
rect 29052 16408 29101 16436
rect 29052 16396 29058 16408
rect 29089 16405 29101 16408
rect 29135 16405 29147 16439
rect 29089 16399 29147 16405
rect 29914 16396 29920 16448
rect 29972 16436 29978 16448
rect 30193 16439 30251 16445
rect 30193 16436 30205 16439
rect 29972 16408 30205 16436
rect 29972 16396 29978 16408
rect 30193 16405 30205 16408
rect 30239 16405 30251 16439
rect 30193 16399 30251 16405
rect 30466 16396 30472 16448
rect 30524 16436 30530 16448
rect 30561 16439 30619 16445
rect 30561 16436 30573 16439
rect 30524 16408 30573 16436
rect 30524 16396 30530 16408
rect 30561 16405 30573 16408
rect 30607 16405 30619 16439
rect 30561 16399 30619 16405
rect 32766 16396 32772 16448
rect 32824 16436 32830 16448
rect 33226 16436 33232 16448
rect 32824 16408 33232 16436
rect 32824 16396 32830 16408
rect 33226 16396 33232 16408
rect 33284 16396 33290 16448
rect 33413 16439 33471 16445
rect 33413 16405 33425 16439
rect 33459 16436 33471 16439
rect 33686 16436 33692 16448
rect 33459 16408 33692 16436
rect 33459 16405 33471 16408
rect 33413 16399 33471 16405
rect 33686 16396 33692 16408
rect 33744 16396 33750 16448
rect 33870 16396 33876 16448
rect 33928 16436 33934 16448
rect 35989 16439 36047 16445
rect 35989 16436 36001 16439
rect 33928 16408 36001 16436
rect 33928 16396 33934 16408
rect 35989 16405 36001 16408
rect 36035 16405 36047 16439
rect 35989 16399 36047 16405
rect 36354 16396 36360 16448
rect 36412 16436 36418 16448
rect 36633 16439 36691 16445
rect 36633 16436 36645 16439
rect 36412 16408 36645 16436
rect 36412 16396 36418 16408
rect 36633 16405 36645 16408
rect 36679 16405 36691 16439
rect 36633 16399 36691 16405
rect 1104 16346 39352 16368
rect 1104 16294 10472 16346
rect 10524 16294 10536 16346
rect 10588 16294 10600 16346
rect 10652 16294 10664 16346
rect 10716 16294 10728 16346
rect 10780 16294 19994 16346
rect 20046 16294 20058 16346
rect 20110 16294 20122 16346
rect 20174 16294 20186 16346
rect 20238 16294 20250 16346
rect 20302 16294 29516 16346
rect 29568 16294 29580 16346
rect 29632 16294 29644 16346
rect 29696 16294 29708 16346
rect 29760 16294 29772 16346
rect 29824 16294 39038 16346
rect 39090 16294 39102 16346
rect 39154 16294 39166 16346
rect 39218 16294 39230 16346
rect 39282 16294 39294 16346
rect 39346 16294 39352 16346
rect 1104 16272 39352 16294
rect 2682 16192 2688 16244
rect 2740 16232 2746 16244
rect 8570 16232 8576 16244
rect 2740 16204 8576 16232
rect 2740 16192 2746 16204
rect 8570 16192 8576 16204
rect 8628 16192 8634 16244
rect 10962 16232 10968 16244
rect 8956 16204 10968 16232
rect 3234 16124 3240 16176
rect 3292 16124 3298 16176
rect 5626 16124 5632 16176
rect 5684 16124 5690 16176
rect 6822 16124 6828 16176
rect 6880 16164 6886 16176
rect 8956 16173 8984 16204
rect 10962 16192 10968 16204
rect 11020 16232 11026 16244
rect 11020 16204 11284 16232
rect 11020 16192 11026 16204
rect 8941 16167 8999 16173
rect 8941 16164 8953 16167
rect 6880 16136 8953 16164
rect 6880 16124 6886 16136
rect 8941 16133 8953 16136
rect 8987 16133 8999 16167
rect 8941 16127 8999 16133
rect 9122 16124 9128 16176
rect 9180 16124 9186 16176
rect 1578 16056 1584 16108
rect 1636 16056 1642 16108
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 5077 16099 5135 16105
rect 5077 16096 5089 16099
rect 4580 16068 5089 16096
rect 4580 16056 4586 16068
rect 5077 16065 5089 16068
rect 5123 16096 5135 16099
rect 5123 16068 8800 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 2222 15988 2228 16040
rect 2280 15988 2286 16040
rect 2498 15988 2504 16040
rect 2556 15988 2562 16040
rect 5166 15988 5172 16040
rect 5224 16028 5230 16040
rect 7742 16028 7748 16040
rect 5224 16000 7748 16028
rect 5224 15988 5230 16000
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 8662 15920 8668 15972
rect 8720 15920 8726 15972
rect 8772 15960 8800 16068
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 10965 16099 11023 16105
rect 10965 16096 10977 16099
rect 9732 16068 10977 16096
rect 9732 16056 9738 16068
rect 10965 16065 10977 16068
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 9214 15988 9220 16040
rect 9272 15988 9278 16040
rect 10980 16028 11008 16059
rect 11256 16028 11284 16204
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 11793 16235 11851 16241
rect 11793 16232 11805 16235
rect 11756 16204 11805 16232
rect 11756 16192 11762 16204
rect 11793 16201 11805 16204
rect 11839 16201 11851 16235
rect 11793 16195 11851 16201
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 21818 16232 21824 16244
rect 12768 16204 21824 16232
rect 12768 16192 12774 16204
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 23198 16232 23204 16244
rect 22296 16204 23204 16232
rect 12437 16167 12495 16173
rect 12437 16133 12449 16167
rect 12483 16164 12495 16167
rect 12618 16164 12624 16176
rect 12483 16136 12624 16164
rect 12483 16133 12495 16136
rect 12437 16127 12495 16133
rect 12618 16124 12624 16136
rect 12676 16124 12682 16176
rect 13538 16124 13544 16176
rect 13596 16124 13602 16176
rect 14182 16124 14188 16176
rect 14240 16124 14246 16176
rect 15102 16124 15108 16176
rect 15160 16164 15166 16176
rect 22296 16173 22324 16204
rect 23198 16192 23204 16204
rect 23256 16192 23262 16244
rect 23566 16192 23572 16244
rect 23624 16232 23630 16244
rect 23753 16235 23811 16241
rect 23753 16232 23765 16235
rect 23624 16204 23765 16232
rect 23624 16192 23630 16204
rect 23753 16201 23765 16204
rect 23799 16201 23811 16235
rect 23753 16195 23811 16201
rect 27522 16192 27528 16244
rect 27580 16192 27586 16244
rect 29178 16192 29184 16244
rect 29236 16192 29242 16244
rect 29840 16204 31248 16232
rect 17129 16167 17187 16173
rect 17129 16164 17141 16167
rect 15160 16136 17141 16164
rect 15160 16124 15166 16136
rect 17129 16133 17141 16136
rect 17175 16133 17187 16167
rect 17129 16127 17187 16133
rect 22281 16167 22339 16173
rect 22281 16133 22293 16167
rect 22327 16133 22339 16167
rect 27540 16164 27568 16192
rect 29840 16164 29868 16204
rect 23506 16136 27568 16164
rect 28934 16136 29868 16164
rect 22281 16127 22339 16133
rect 29914 16124 29920 16176
rect 29972 16124 29978 16176
rect 30926 16124 30932 16176
rect 30984 16124 30990 16176
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16096 11759 16099
rect 11790 16096 11796 16108
rect 11747 16068 11796 16096
rect 11747 16065 11759 16068
rect 11701 16059 11759 16065
rect 11790 16056 11796 16068
rect 11848 16056 11854 16108
rect 13170 16056 13176 16108
rect 13228 16096 13234 16108
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 13228 16068 13277 16096
rect 13228 16056 13234 16068
rect 13265 16065 13277 16068
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 15378 16056 15384 16108
rect 15436 16096 15442 16108
rect 15841 16099 15899 16105
rect 15841 16096 15853 16099
rect 15436 16068 15853 16096
rect 15436 16056 15442 16068
rect 15841 16065 15853 16068
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 16022 16056 16028 16108
rect 16080 16056 16086 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16390 16096 16396 16108
rect 16163 16068 16396 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16096 16911 16099
rect 20346 16096 20352 16108
rect 16899 16068 20352 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 20346 16056 20352 16068
rect 20404 16056 20410 16108
rect 27338 16056 27344 16108
rect 27396 16096 27402 16108
rect 27433 16099 27491 16105
rect 27433 16096 27445 16099
rect 27396 16068 27445 16096
rect 27396 16056 27402 16068
rect 27433 16065 27445 16068
rect 27479 16065 27491 16099
rect 27433 16059 27491 16065
rect 10980 16000 11192 16028
rect 11256 16000 14964 16028
rect 8772 15932 10180 15960
rect 1673 15895 1731 15901
rect 1673 15861 1685 15895
rect 1719 15892 1731 15895
rect 2958 15892 2964 15904
rect 1719 15864 2964 15892
rect 1719 15861 1731 15864
rect 1673 15855 1731 15861
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 3142 15852 3148 15904
rect 3200 15892 3206 15904
rect 3973 15895 4031 15901
rect 3973 15892 3985 15895
rect 3200 15864 3985 15892
rect 3200 15852 3206 15864
rect 3973 15861 3985 15864
rect 4019 15892 4031 15895
rect 10042 15892 10048 15904
rect 4019 15864 10048 15892
rect 4019 15861 4031 15864
rect 3973 15855 4031 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 10152 15892 10180 15932
rect 11054 15920 11060 15972
rect 11112 15920 11118 15972
rect 11164 15960 11192 16000
rect 11164 15932 12664 15960
rect 11882 15892 11888 15904
rect 10152 15864 11888 15892
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 12636 15892 12664 15932
rect 12710 15920 12716 15972
rect 12768 15960 12774 15972
rect 12894 15960 12900 15972
rect 12768 15932 12900 15960
rect 12768 15920 12774 15932
rect 12894 15920 12900 15932
rect 12952 15920 12958 15972
rect 13998 15892 14004 15904
rect 12636 15864 14004 15892
rect 13998 15852 14004 15864
rect 14056 15852 14062 15904
rect 14936 15892 14964 16000
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 15746 15988 15752 16040
rect 15804 16028 15810 16040
rect 16298 16028 16304 16040
rect 15804 16000 16304 16028
rect 15804 15988 15810 16000
rect 16298 15988 16304 16000
rect 16356 15988 16362 16040
rect 20714 15988 20720 16040
rect 20772 16028 20778 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 20772 16000 22017 16028
rect 20772 15988 20778 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 22370 15988 22376 16040
rect 22428 16028 22434 16040
rect 26694 16028 26700 16040
rect 22428 16000 26700 16028
rect 22428 15988 22434 16000
rect 26694 15988 26700 16000
rect 26752 15988 26758 16040
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 16028 27767 16031
rect 29362 16028 29368 16040
rect 27755 16000 29368 16028
rect 27755 15997 27767 16000
rect 27709 15991 27767 15997
rect 29362 15988 29368 16000
rect 29420 15988 29426 16040
rect 29641 16031 29699 16037
rect 29641 15997 29653 16031
rect 29687 16028 29699 16031
rect 31220 16028 31248 16204
rect 33686 16192 33692 16244
rect 33744 16232 33750 16244
rect 35342 16232 35348 16244
rect 33744 16204 35348 16232
rect 33744 16192 33750 16204
rect 35342 16192 35348 16204
rect 35400 16192 35406 16244
rect 33042 16164 33048 16176
rect 32508 16136 33048 16164
rect 31294 16056 31300 16108
rect 31352 16096 31358 16108
rect 32508 16105 32536 16136
rect 33042 16124 33048 16136
rect 33100 16124 33106 16176
rect 33318 16124 33324 16176
rect 33376 16164 33382 16176
rect 33413 16167 33471 16173
rect 33413 16164 33425 16167
rect 33376 16136 33425 16164
rect 33376 16124 33382 16136
rect 33413 16133 33425 16136
rect 33459 16133 33471 16167
rect 34698 16164 34704 16176
rect 34638 16136 34704 16164
rect 33413 16127 33471 16133
rect 34698 16124 34704 16136
rect 34756 16124 34762 16176
rect 35066 16124 35072 16176
rect 35124 16164 35130 16176
rect 38470 16164 38476 16176
rect 35124 16136 38476 16164
rect 35124 16124 35130 16136
rect 38470 16124 38476 16136
rect 38528 16124 38534 16176
rect 32493 16099 32551 16105
rect 32493 16096 32505 16099
rect 31352 16068 32505 16096
rect 31352 16056 31358 16068
rect 32493 16065 32505 16068
rect 32539 16065 32551 16099
rect 32493 16059 32551 16065
rect 32950 16056 32956 16108
rect 33008 16096 33014 16108
rect 33137 16099 33195 16105
rect 33137 16096 33149 16099
rect 33008 16068 33149 16096
rect 33008 16056 33014 16068
rect 33137 16065 33149 16068
rect 33183 16065 33195 16099
rect 33137 16059 33195 16065
rect 35802 16056 35808 16108
rect 35860 16096 35866 16108
rect 35860 16068 36584 16096
rect 35860 16056 35866 16068
rect 33870 16028 33876 16040
rect 29687 16000 29776 16028
rect 31220 16000 33876 16028
rect 29687 15997 29699 16000
rect 29641 15991 29699 15997
rect 15194 15920 15200 15972
rect 15252 15960 15258 15972
rect 15565 15963 15623 15969
rect 15565 15960 15577 15963
rect 15252 15932 15577 15960
rect 15252 15920 15258 15932
rect 15565 15929 15577 15932
rect 15611 15929 15623 15963
rect 15565 15923 15623 15929
rect 15933 15963 15991 15969
rect 15933 15929 15945 15963
rect 15979 15960 15991 15963
rect 17862 15960 17868 15972
rect 15979 15932 17868 15960
rect 15979 15929 15991 15932
rect 15933 15923 15991 15929
rect 17862 15920 17868 15932
rect 17920 15920 17926 15972
rect 19886 15892 19892 15904
rect 14936 15864 19892 15892
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 22738 15852 22744 15904
rect 22796 15892 22802 15904
rect 28718 15892 28724 15904
rect 22796 15864 28724 15892
rect 22796 15852 22802 15864
rect 28718 15852 28724 15864
rect 28776 15852 28782 15904
rect 29748 15892 29776 16000
rect 33870 15988 33876 16000
rect 33928 15988 33934 16040
rect 34146 15988 34152 16040
rect 34204 16028 34210 16040
rect 35897 16031 35955 16037
rect 35897 16028 35909 16031
rect 34204 16000 35909 16028
rect 34204 15988 34210 16000
rect 35897 15997 35909 16000
rect 35943 15997 35955 16031
rect 35897 15991 35955 15997
rect 35989 16031 36047 16037
rect 35989 15997 36001 16031
rect 36035 15997 36047 16031
rect 36556 16028 36584 16068
rect 36630 16056 36636 16108
rect 36688 16096 36694 16108
rect 37182 16096 37188 16108
rect 36688 16068 37188 16096
rect 36688 16056 36694 16068
rect 37182 16056 37188 16068
rect 37240 16056 37246 16108
rect 37461 16099 37519 16105
rect 37461 16065 37473 16099
rect 37507 16096 37519 16099
rect 37550 16096 37556 16108
rect 37507 16068 37556 16096
rect 37507 16065 37519 16068
rect 37461 16059 37519 16065
rect 37550 16056 37556 16068
rect 37608 16056 37614 16108
rect 37918 16028 37924 16040
rect 36556 16000 37924 16028
rect 35989 15991 36047 15997
rect 30926 15920 30932 15972
rect 30984 15960 30990 15972
rect 30984 15932 32720 15960
rect 30984 15920 30990 15932
rect 30282 15892 30288 15904
rect 29748 15864 30288 15892
rect 30282 15852 30288 15864
rect 30340 15852 30346 15904
rect 30650 15852 30656 15904
rect 30708 15892 30714 15904
rect 31389 15895 31447 15901
rect 31389 15892 31401 15895
rect 30708 15864 31401 15892
rect 30708 15852 30714 15864
rect 31389 15861 31401 15864
rect 31435 15861 31447 15895
rect 31389 15855 31447 15861
rect 32582 15852 32588 15904
rect 32640 15852 32646 15904
rect 32692 15892 32720 15932
rect 34790 15920 34796 15972
rect 34848 15960 34854 15972
rect 36004 15960 36032 15991
rect 37918 15988 37924 16000
rect 37976 15988 37982 16040
rect 34848 15932 36032 15960
rect 34848 15920 34854 15932
rect 34146 15892 34152 15904
rect 32692 15864 34152 15892
rect 34146 15852 34152 15864
rect 34204 15852 34210 15904
rect 34882 15852 34888 15904
rect 34940 15852 34946 15904
rect 35434 15852 35440 15904
rect 35492 15852 35498 15904
rect 36722 15852 36728 15904
rect 36780 15852 36786 15904
rect 37274 15852 37280 15904
rect 37332 15892 37338 15904
rect 37553 15895 37611 15901
rect 37553 15892 37565 15895
rect 37332 15864 37565 15892
rect 37332 15852 37338 15864
rect 37553 15861 37565 15864
rect 37599 15861 37611 15895
rect 37553 15855 37611 15861
rect 1104 15802 39192 15824
rect 1104 15750 5711 15802
rect 5763 15750 5775 15802
rect 5827 15750 5839 15802
rect 5891 15750 5903 15802
rect 5955 15750 5967 15802
rect 6019 15750 15233 15802
rect 15285 15750 15297 15802
rect 15349 15750 15361 15802
rect 15413 15750 15425 15802
rect 15477 15750 15489 15802
rect 15541 15750 24755 15802
rect 24807 15750 24819 15802
rect 24871 15750 24883 15802
rect 24935 15750 24947 15802
rect 24999 15750 25011 15802
rect 25063 15750 34277 15802
rect 34329 15750 34341 15802
rect 34393 15750 34405 15802
rect 34457 15750 34469 15802
rect 34521 15750 34533 15802
rect 34585 15750 39192 15802
rect 1104 15728 39192 15750
rect 2498 15648 2504 15700
rect 2556 15688 2562 15700
rect 2685 15691 2743 15697
rect 2685 15688 2697 15691
rect 2556 15660 2697 15688
rect 2556 15648 2562 15660
rect 2685 15657 2697 15660
rect 2731 15657 2743 15691
rect 2685 15651 2743 15657
rect 3602 15648 3608 15700
rect 3660 15688 3666 15700
rect 5721 15691 5779 15697
rect 5721 15688 5733 15691
rect 3660 15660 5733 15688
rect 3660 15648 3666 15660
rect 5721 15657 5733 15660
rect 5767 15657 5779 15691
rect 5721 15651 5779 15657
rect 5828 15660 7052 15688
rect 3142 15512 3148 15564
rect 3200 15512 3206 15564
rect 3326 15512 3332 15564
rect 3384 15512 3390 15564
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 5828 15552 5856 15660
rect 4672 15524 5856 15552
rect 7024 15552 7052 15660
rect 8202 15648 8208 15700
rect 8260 15648 8266 15700
rect 10032 15691 10090 15697
rect 10032 15657 10044 15691
rect 10078 15688 10090 15691
rect 11698 15688 11704 15700
rect 10078 15660 11704 15688
rect 10078 15657 10090 15660
rect 10032 15651 10090 15657
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 13630 15688 13636 15700
rect 11940 15660 13636 15688
rect 11940 15648 11946 15660
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 13722 15648 13728 15700
rect 13780 15648 13786 15700
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 15102 15688 15108 15700
rect 14240 15660 15108 15688
rect 14240 15648 14246 15660
rect 15102 15648 15108 15660
rect 15160 15648 15166 15700
rect 15212 15660 26372 15688
rect 15212 15620 15240 15660
rect 13244 15592 15240 15620
rect 19797 15623 19855 15629
rect 9217 15555 9275 15561
rect 9217 15552 9229 15555
rect 7024 15524 9229 15552
rect 4672 15512 4678 15524
rect 9217 15521 9229 15524
rect 9263 15521 9275 15555
rect 9217 15515 9275 15521
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 11977 15555 12035 15561
rect 11977 15552 11989 15555
rect 9824 15524 11989 15552
rect 9824 15512 9830 15524
rect 11977 15521 11989 15524
rect 12023 15552 12035 15555
rect 12618 15552 12624 15564
rect 12023 15524 12624 15552
rect 12023 15521 12035 15524
rect 11977 15515 12035 15521
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 13244 15552 13272 15592
rect 19797 15589 19809 15623
rect 19843 15620 19855 15623
rect 19978 15620 19984 15632
rect 19843 15592 19984 15620
rect 19843 15589 19855 15592
rect 19797 15583 19855 15589
rect 19978 15580 19984 15592
rect 20036 15620 20042 15632
rect 20622 15620 20628 15632
rect 20036 15592 20628 15620
rect 20036 15580 20042 15592
rect 20622 15580 20628 15592
rect 20680 15580 20686 15632
rect 24854 15580 24860 15632
rect 24912 15620 24918 15632
rect 25225 15623 25283 15629
rect 25225 15620 25237 15623
rect 24912 15592 25237 15620
rect 24912 15580 24918 15592
rect 25225 15589 25237 15592
rect 25271 15589 25283 15623
rect 26344 15620 26372 15660
rect 26418 15648 26424 15700
rect 26476 15648 26482 15700
rect 27614 15648 27620 15700
rect 27672 15688 27678 15700
rect 28445 15691 28503 15697
rect 28445 15688 28457 15691
rect 27672 15660 28457 15688
rect 27672 15648 27678 15660
rect 28445 15657 28457 15660
rect 28491 15657 28503 15691
rect 28445 15651 28503 15657
rect 28718 15648 28724 15700
rect 28776 15688 28782 15700
rect 30926 15688 30932 15700
rect 28776 15660 30932 15688
rect 28776 15648 28782 15660
rect 30926 15648 30932 15660
rect 30984 15648 30990 15700
rect 31202 15648 31208 15700
rect 31260 15688 31266 15700
rect 33873 15691 33931 15697
rect 33873 15688 33885 15691
rect 31260 15660 33885 15688
rect 31260 15648 31266 15660
rect 33873 15657 33885 15660
rect 33919 15657 33931 15691
rect 33873 15651 33931 15657
rect 34057 15691 34115 15697
rect 34057 15657 34069 15691
rect 34103 15688 34115 15691
rect 35986 15688 35992 15700
rect 34103 15660 35992 15688
rect 34103 15657 34115 15660
rect 34057 15651 34115 15657
rect 35986 15648 35992 15660
rect 36044 15648 36050 15700
rect 28077 15623 28135 15629
rect 28077 15620 28089 15623
rect 26344 15592 28089 15620
rect 25225 15583 25283 15589
rect 28077 15589 28089 15592
rect 28123 15589 28135 15623
rect 28077 15583 28135 15589
rect 12952 15524 13272 15552
rect 12952 15512 12958 15524
rect 14090 15512 14096 15564
rect 14148 15552 14154 15564
rect 15933 15555 15991 15561
rect 15933 15552 15945 15555
rect 14148 15524 15945 15552
rect 14148 15512 14154 15524
rect 15933 15521 15945 15524
rect 15979 15521 15991 15555
rect 15933 15515 15991 15521
rect 16209 15555 16267 15561
rect 16209 15521 16221 15555
rect 16255 15552 16267 15555
rect 16850 15552 16856 15564
rect 16255 15524 16856 15552
rect 16255 15521 16267 15524
rect 16209 15515 16267 15521
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 22833 15555 22891 15561
rect 22833 15521 22845 15555
rect 22879 15552 22891 15555
rect 25685 15555 25743 15561
rect 22879 15524 25636 15552
rect 22879 15521 22891 15524
rect 22833 15515 22891 15521
rect 934 15444 940 15496
rect 992 15484 998 15496
rect 1581 15487 1639 15493
rect 1581 15484 1593 15487
rect 992 15456 1593 15484
rect 992 15444 998 15456
rect 1581 15453 1593 15456
rect 1627 15453 1639 15487
rect 1581 15447 1639 15453
rect 3970 15444 3976 15496
rect 4028 15444 4034 15496
rect 5626 15444 5632 15496
rect 5684 15484 5690 15496
rect 6181 15487 6239 15493
rect 6181 15484 6193 15487
rect 5684 15456 6193 15484
rect 5684 15444 5690 15456
rect 6181 15453 6193 15456
rect 6227 15453 6239 15487
rect 6181 15447 6239 15453
rect 6638 15444 6644 15496
rect 6696 15484 6702 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6696 15456 6837 15484
rect 6696 15444 6702 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 7558 15444 7564 15496
rect 7616 15484 7622 15496
rect 8113 15487 8171 15493
rect 8113 15484 8125 15487
rect 7616 15456 8125 15484
rect 7616 15444 7622 15456
rect 8113 15453 8125 15456
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9674 15484 9680 15496
rect 9171 15456 9680 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 14366 15484 14372 15496
rect 13386 15456 14372 15484
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 17954 15484 17960 15496
rect 17342 15456 17960 15484
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15484 19579 15487
rect 20346 15484 20352 15496
rect 19567 15456 20352 15484
rect 19567 15453 19579 15456
rect 19521 15447 19579 15453
rect 1857 15419 1915 15425
rect 1857 15385 1869 15419
rect 1903 15416 1915 15419
rect 2682 15416 2688 15428
rect 1903 15388 2688 15416
rect 1903 15385 1915 15388
rect 1857 15379 1915 15385
rect 2682 15376 2688 15388
rect 2740 15376 2746 15428
rect 4154 15376 4160 15428
rect 4212 15416 4218 15428
rect 4249 15419 4307 15425
rect 4249 15416 4261 15419
rect 4212 15388 4261 15416
rect 4212 15376 4218 15388
rect 4249 15385 4261 15388
rect 4295 15385 4307 15419
rect 4249 15379 4307 15385
rect 4706 15376 4712 15428
rect 4764 15376 4770 15428
rect 6273 15419 6331 15425
rect 6273 15385 6285 15419
rect 6319 15416 6331 15419
rect 12253 15419 12311 15425
rect 6319 15388 10534 15416
rect 6319 15385 6331 15388
rect 6273 15379 6331 15385
rect 12253 15385 12265 15419
rect 12299 15416 12311 15419
rect 12342 15416 12348 15428
rect 12299 15388 12348 15416
rect 12299 15385 12311 15388
rect 12253 15379 12311 15385
rect 12342 15376 12348 15388
rect 12400 15376 12406 15428
rect 14274 15376 14280 15428
rect 14332 15376 14338 15428
rect 15010 15416 15016 15428
rect 14384 15388 15016 15416
rect 3050 15308 3056 15360
rect 3108 15308 3114 15360
rect 6917 15351 6975 15357
rect 6917 15317 6929 15351
rect 6963 15348 6975 15351
rect 8202 15348 8208 15360
rect 6963 15320 8208 15348
rect 6963 15317 6975 15320
rect 6917 15311 6975 15317
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 10134 15348 10140 15360
rect 8352 15320 10140 15348
rect 8352 15308 8358 15320
rect 10134 15308 10140 15320
rect 10192 15308 10198 15360
rect 11517 15351 11575 15357
rect 11517 15317 11529 15351
rect 11563 15348 11575 15351
rect 11882 15348 11888 15360
rect 11563 15320 11888 15348
rect 11563 15317 11575 15320
rect 11517 15311 11575 15317
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 14384 15348 14412 15388
rect 15010 15376 15016 15388
rect 15068 15376 15074 15428
rect 18156 15416 18184 15447
rect 20346 15444 20352 15456
rect 20404 15444 20410 15496
rect 20714 15444 20720 15496
rect 20772 15484 20778 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 20772 15456 21097 15484
rect 20772 15444 20778 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 23842 15444 23848 15496
rect 23900 15444 23906 15496
rect 25608 15484 25636 15524
rect 25685 15521 25697 15555
rect 25731 15552 25743 15555
rect 26602 15552 26608 15564
rect 25731 15524 26608 15552
rect 25731 15521 25743 15524
rect 25685 15515 25743 15521
rect 26602 15512 26608 15524
rect 26660 15512 26666 15564
rect 26234 15484 26240 15496
rect 25608 15456 26240 15484
rect 26234 15444 26240 15456
rect 26292 15444 26298 15496
rect 26326 15444 26332 15496
rect 26384 15444 26390 15496
rect 28092 15484 28120 15583
rect 28166 15580 28172 15632
rect 28224 15620 28230 15632
rect 28534 15620 28540 15632
rect 28224 15592 28540 15620
rect 28224 15580 28230 15592
rect 28534 15580 28540 15592
rect 28592 15620 28598 15632
rect 31294 15620 31300 15632
rect 28592 15592 29040 15620
rect 28592 15580 28598 15592
rect 28902 15512 28908 15564
rect 28960 15512 28966 15564
rect 29012 15561 29040 15592
rect 30208 15592 31300 15620
rect 30208 15564 30236 15592
rect 31294 15580 31300 15592
rect 31352 15580 31358 15632
rect 31754 15580 31760 15632
rect 31812 15620 31818 15632
rect 32769 15623 32827 15629
rect 32769 15620 32781 15623
rect 31812 15592 32781 15620
rect 31812 15580 31818 15592
rect 32769 15589 32781 15592
rect 32815 15589 32827 15623
rect 32769 15583 32827 15589
rect 32861 15623 32919 15629
rect 32861 15589 32873 15623
rect 32907 15620 32919 15623
rect 32950 15620 32956 15632
rect 32907 15592 32956 15620
rect 32907 15589 32919 15592
rect 32861 15583 32919 15589
rect 32950 15580 32956 15592
rect 33008 15580 33014 15632
rect 34900 15592 35204 15620
rect 28997 15555 29055 15561
rect 28997 15521 29009 15555
rect 29043 15521 29055 15555
rect 28997 15515 29055 15521
rect 30190 15512 30196 15564
rect 30248 15512 30254 15564
rect 33778 15552 33784 15564
rect 33060 15524 33784 15552
rect 28813 15487 28871 15493
rect 28813 15484 28825 15487
rect 28092 15456 28825 15484
rect 28813 15453 28825 15456
rect 28859 15453 28871 15487
rect 28813 15447 28871 15453
rect 29914 15444 29920 15496
rect 29972 15444 29978 15496
rect 31386 15444 31392 15496
rect 31444 15444 31450 15496
rect 31478 15444 31484 15496
rect 31536 15484 31542 15496
rect 31665 15487 31723 15493
rect 31665 15484 31677 15487
rect 31536 15456 31677 15484
rect 31536 15444 31542 15456
rect 31665 15453 31677 15456
rect 31711 15453 31723 15487
rect 31665 15447 31723 15453
rect 31757 15487 31815 15493
rect 31757 15453 31769 15487
rect 31803 15484 31815 15487
rect 31803 15456 31892 15484
rect 31803 15453 31815 15456
rect 31757 15447 31815 15453
rect 19150 15416 19156 15428
rect 17604 15388 19156 15416
rect 12676 15320 14412 15348
rect 12676 15308 12682 15320
rect 14826 15308 14832 15360
rect 14884 15348 14890 15360
rect 17604 15348 17632 15388
rect 19150 15376 19156 15388
rect 19208 15416 19214 15428
rect 19702 15416 19708 15428
rect 19208 15388 19708 15416
rect 19208 15376 19214 15388
rect 19702 15376 19708 15388
rect 19760 15376 19766 15428
rect 20070 15376 20076 15428
rect 20128 15416 20134 15428
rect 20898 15416 20904 15428
rect 20128 15388 20904 15416
rect 20128 15376 20134 15388
rect 20898 15376 20904 15388
rect 20956 15376 20962 15428
rect 21361 15419 21419 15425
rect 21361 15385 21373 15419
rect 21407 15385 21419 15419
rect 21361 15379 21419 15385
rect 14884 15320 17632 15348
rect 14884 15308 14890 15320
rect 17678 15308 17684 15360
rect 17736 15308 17742 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18325 15351 18383 15357
rect 18325 15348 18337 15351
rect 18012 15320 18337 15348
rect 18012 15308 18018 15320
rect 18325 15317 18337 15320
rect 18371 15348 18383 15351
rect 19426 15348 19432 15360
rect 18371 15320 19432 15348
rect 18371 15317 18383 15320
rect 18325 15311 18383 15317
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 21376 15348 21404 15379
rect 21818 15376 21824 15428
rect 21876 15376 21882 15428
rect 25498 15416 25504 15428
rect 22756 15388 25504 15416
rect 22756 15348 22784 15388
rect 25498 15376 25504 15388
rect 25556 15376 25562 15428
rect 25774 15376 25780 15428
rect 25832 15376 25838 15428
rect 26694 15376 26700 15428
rect 26752 15416 26758 15428
rect 31570 15416 31576 15428
rect 26752 15388 31576 15416
rect 26752 15376 26758 15388
rect 31570 15376 31576 15388
rect 31628 15376 31634 15428
rect 21376 15320 22784 15348
rect 23934 15308 23940 15360
rect 23992 15308 23998 15360
rect 24857 15351 24915 15357
rect 24857 15317 24869 15351
rect 24903 15348 24915 15351
rect 25682 15348 25688 15360
rect 24903 15320 25688 15348
rect 24903 15317 24915 15320
rect 24857 15311 24915 15317
rect 25682 15308 25688 15320
rect 25740 15308 25746 15360
rect 28810 15308 28816 15360
rect 28868 15348 28874 15360
rect 31110 15348 31116 15360
rect 28868 15320 31116 15348
rect 28868 15308 28874 15320
rect 31110 15308 31116 15320
rect 31168 15348 31174 15360
rect 31864 15348 31892 15456
rect 32214 15444 32220 15496
rect 32272 15484 32278 15496
rect 33060 15493 33088 15524
rect 33778 15512 33784 15524
rect 33836 15512 33842 15564
rect 32953 15487 33011 15493
rect 32953 15484 32965 15487
rect 32272 15456 32965 15484
rect 32272 15444 32278 15456
rect 32953 15453 32965 15456
rect 32999 15453 33011 15487
rect 32953 15447 33011 15453
rect 33045 15487 33103 15493
rect 33045 15453 33057 15487
rect 33091 15453 33103 15487
rect 33045 15447 33103 15453
rect 33226 15444 33232 15496
rect 33284 15484 33290 15496
rect 33502 15484 33508 15496
rect 33284 15456 33508 15484
rect 33284 15444 33290 15456
rect 33502 15444 33508 15456
rect 33560 15444 33566 15496
rect 34900 15484 34928 15592
rect 35066 15512 35072 15564
rect 35124 15512 35130 15564
rect 35176 15552 35204 15592
rect 36446 15580 36452 15632
rect 36504 15620 36510 15632
rect 36504 15592 38148 15620
rect 36504 15580 36510 15592
rect 37366 15552 37372 15564
rect 35176 15524 37372 15552
rect 37366 15512 37372 15524
rect 37424 15512 37430 15564
rect 38120 15561 38148 15592
rect 38105 15555 38163 15561
rect 38105 15521 38117 15555
rect 38151 15521 38163 15555
rect 38105 15515 38163 15521
rect 33612 15456 34928 15484
rect 32493 15419 32551 15425
rect 32493 15385 32505 15419
rect 32539 15416 32551 15419
rect 33612 15416 33640 15456
rect 37918 15444 37924 15496
rect 37976 15444 37982 15496
rect 32539 15388 33640 15416
rect 33689 15419 33747 15425
rect 32539 15385 32551 15388
rect 32493 15379 32551 15385
rect 33689 15385 33701 15419
rect 33735 15416 33747 15419
rect 34146 15416 34152 15428
rect 33735 15388 34152 15416
rect 33735 15385 33747 15388
rect 33689 15379 33747 15385
rect 34146 15376 34152 15388
rect 34204 15376 34210 15428
rect 35345 15419 35403 15425
rect 35345 15385 35357 15419
rect 35391 15385 35403 15419
rect 36722 15416 36728 15428
rect 36570 15388 36728 15416
rect 35345 15379 35403 15385
rect 31168 15320 31892 15348
rect 31941 15351 31999 15357
rect 31168 15308 31174 15320
rect 31941 15317 31953 15351
rect 31987 15348 31999 15351
rect 32030 15348 32036 15360
rect 31987 15320 32036 15348
rect 31987 15317 31999 15320
rect 31941 15311 31999 15317
rect 32030 15308 32036 15320
rect 32088 15308 32094 15360
rect 32122 15308 32128 15360
rect 32180 15348 32186 15360
rect 33226 15348 33232 15360
rect 32180 15320 33232 15348
rect 32180 15308 32186 15320
rect 33226 15308 33232 15320
rect 33284 15308 33290 15360
rect 33410 15308 33416 15360
rect 33468 15348 33474 15360
rect 33889 15351 33947 15357
rect 33889 15348 33901 15351
rect 33468 15320 33901 15348
rect 33468 15308 33474 15320
rect 33889 15317 33901 15320
rect 33935 15317 33947 15351
rect 35360 15348 35388 15379
rect 36722 15376 36728 15388
rect 36780 15376 36786 15428
rect 37090 15376 37096 15428
rect 37148 15416 37154 15428
rect 38013 15419 38071 15425
rect 38013 15416 38025 15419
rect 37148 15388 38025 15416
rect 37148 15376 37154 15388
rect 38013 15385 38025 15388
rect 38059 15385 38071 15419
rect 38013 15379 38071 15385
rect 37553 15351 37611 15357
rect 37553 15348 37565 15351
rect 35360 15320 37565 15348
rect 33889 15311 33947 15317
rect 37553 15317 37565 15320
rect 37599 15317 37611 15351
rect 37553 15311 37611 15317
rect 1104 15258 39352 15280
rect 1104 15206 10472 15258
rect 10524 15206 10536 15258
rect 10588 15206 10600 15258
rect 10652 15206 10664 15258
rect 10716 15206 10728 15258
rect 10780 15206 19994 15258
rect 20046 15206 20058 15258
rect 20110 15206 20122 15258
rect 20174 15206 20186 15258
rect 20238 15206 20250 15258
rect 20302 15206 29516 15258
rect 29568 15206 29580 15258
rect 29632 15206 29644 15258
rect 29696 15206 29708 15258
rect 29760 15206 29772 15258
rect 29824 15206 39038 15258
rect 39090 15206 39102 15258
rect 39154 15206 39166 15258
rect 39218 15206 39230 15258
rect 39282 15206 39294 15258
rect 39346 15206 39352 15258
rect 1104 15184 39352 15206
rect 4890 15144 4896 15156
rect 2240 15116 4896 15144
rect 2240 15017 2268 15116
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 4982 15104 4988 15156
rect 5040 15144 5046 15156
rect 7101 15147 7159 15153
rect 5040 15116 6500 15144
rect 5040 15104 5046 15116
rect 2590 15036 2596 15088
rect 2648 15076 2654 15088
rect 3237 15079 3295 15085
rect 3237 15076 3249 15079
rect 2648 15048 3249 15076
rect 2648 15036 2654 15048
rect 3237 15045 3249 15048
rect 3283 15045 3295 15079
rect 3237 15039 3295 15045
rect 4246 15036 4252 15088
rect 4304 15036 4310 15088
rect 5534 15036 5540 15088
rect 5592 15036 5598 15088
rect 5626 15036 5632 15088
rect 5684 15076 5690 15088
rect 5721 15079 5779 15085
rect 5721 15076 5733 15079
rect 5684 15048 5733 15076
rect 5684 15036 5690 15048
rect 5721 15045 5733 15048
rect 5767 15045 5779 15079
rect 5721 15039 5779 15045
rect 5813 15079 5871 15085
rect 5813 15045 5825 15079
rect 5859 15076 5871 15079
rect 6362 15076 6368 15088
rect 5859 15048 6368 15076
rect 5859 15045 5871 15048
rect 5813 15039 5871 15045
rect 6362 15036 6368 15048
rect 6420 15036 6426 15088
rect 6472 15076 6500 15116
rect 7101 15113 7113 15147
rect 7147 15144 7159 15147
rect 7147 15116 7604 15144
rect 7147 15113 7159 15116
rect 7101 15107 7159 15113
rect 6825 15079 6883 15085
rect 6825 15076 6837 15079
rect 6472 15048 6837 15076
rect 6825 15045 6837 15048
rect 6871 15045 6883 15079
rect 6825 15039 6883 15045
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 14977 2283 15011
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 2225 14971 2283 14977
rect 5736 14980 6561 15008
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 2314 14940 2320 14952
rect 2087 14912 2320 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 2961 14943 3019 14949
rect 2961 14909 2973 14943
rect 3007 14940 3019 14943
rect 3970 14940 3976 14952
rect 3007 14912 3976 14940
rect 3007 14909 3019 14912
rect 2961 14903 3019 14909
rect 2222 14832 2228 14884
rect 2280 14872 2286 14884
rect 2976 14872 3004 14903
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 2280 14844 3004 14872
rect 2280 14832 2286 14844
rect 5258 14832 5264 14884
rect 5316 14832 5322 14884
rect 5350 14832 5356 14884
rect 5408 14872 5414 14884
rect 5736 14872 5764 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 6730 14968 6736 15020
rect 6788 14968 6794 15020
rect 7576 15017 7604 15116
rect 7926 15104 7932 15156
rect 7984 15104 7990 15156
rect 10318 15104 10324 15156
rect 10376 15104 10382 15156
rect 11057 15147 11115 15153
rect 11057 15113 11069 15147
rect 11103 15144 11115 15147
rect 11238 15144 11244 15156
rect 11103 15116 11244 15144
rect 11103 15113 11115 15116
rect 11057 15107 11115 15113
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 11698 15104 11704 15156
rect 11756 15104 11762 15156
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 11940 15116 12173 15144
rect 11940 15104 11946 15116
rect 12161 15113 12173 15116
rect 12207 15144 12219 15147
rect 12250 15144 12256 15156
rect 12207 15116 12256 15144
rect 12207 15113 12219 15116
rect 12161 15107 12219 15113
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 17405 15147 17463 15153
rect 17405 15144 17417 15147
rect 12406 15116 17417 15144
rect 11146 15076 11152 15088
rect 10074 15048 11152 15076
rect 11146 15036 11152 15048
rect 11204 15036 11210 15088
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 11974 15076 11980 15088
rect 11480 15048 11980 15076
rect 11480 15036 11486 15048
rect 11974 15036 11980 15048
rect 12032 15076 12038 15088
rect 12406 15076 12434 15116
rect 17405 15113 17417 15116
rect 17451 15113 17463 15147
rect 17405 15107 17463 15113
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 18141 15147 18199 15153
rect 18141 15144 18153 15147
rect 18104 15116 18153 15144
rect 18104 15104 18110 15116
rect 18141 15113 18153 15116
rect 18187 15113 18199 15147
rect 18141 15107 18199 15113
rect 18230 15104 18236 15156
rect 18288 15144 18294 15156
rect 18506 15144 18512 15156
rect 18288 15116 18512 15144
rect 18288 15104 18294 15116
rect 18506 15104 18512 15116
rect 18564 15104 18570 15156
rect 21082 15104 21088 15156
rect 21140 15104 21146 15156
rect 22020 15116 22140 15144
rect 12032 15048 12434 15076
rect 13357 15079 13415 15085
rect 12032 15036 12038 15048
rect 13357 15045 13369 15079
rect 13403 15045 13415 15079
rect 13357 15039 13415 15045
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 14977 6975 15011
rect 6917 14971 6975 14977
rect 7561 15011 7619 15017
rect 7561 14977 7573 15011
rect 7607 14977 7619 15011
rect 7561 14971 7619 14977
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 15008 7803 15011
rect 8386 15008 8392 15020
rect 7791 14980 8392 15008
rect 7791 14977 7803 14980
rect 7745 14971 7803 14977
rect 6932 14940 6960 14971
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 10965 15011 11023 15017
rect 10965 14977 10977 15011
rect 11011 15008 11023 15011
rect 11790 15008 11796 15020
rect 11011 14980 11796 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 12066 14968 12072 15020
rect 12124 14968 12130 15020
rect 8110 14940 8116 14952
rect 6932 14912 8116 14940
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 8573 14943 8631 14949
rect 8573 14940 8585 14943
rect 8352 14912 8585 14940
rect 8352 14900 8358 14912
rect 8573 14909 8585 14912
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14940 8907 14943
rect 9858 14940 9864 14952
rect 8895 14912 9864 14940
rect 8895 14909 8907 14912
rect 8849 14903 8907 14909
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 12253 14943 12311 14949
rect 12253 14940 12265 14943
rect 11572 14912 12265 14940
rect 11572 14900 11578 14912
rect 12253 14909 12265 14912
rect 12299 14940 12311 14943
rect 12342 14940 12348 14952
rect 12299 14912 12348 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 13372 14940 13400 15039
rect 14090 15036 14096 15088
rect 14148 15036 14154 15088
rect 16666 15036 16672 15088
rect 16724 15076 16730 15088
rect 16945 15079 17003 15085
rect 16945 15076 16957 15079
rect 16724 15048 16957 15076
rect 16724 15036 16730 15048
rect 16945 15045 16957 15048
rect 16991 15045 17003 15079
rect 16945 15039 17003 15045
rect 17494 15036 17500 15088
rect 17552 15036 17558 15088
rect 18601 15079 18659 15085
rect 18601 15045 18613 15079
rect 18647 15045 18659 15079
rect 18601 15039 18659 15045
rect 13722 14968 13728 15020
rect 13780 15008 13786 15020
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 13780 14980 15485 15008
rect 13780 14968 13786 14980
rect 15473 14977 15485 14980
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 14366 14940 14372 14952
rect 12768 14912 14372 14940
rect 12768 14900 12774 14912
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 15488 14940 15516 14971
rect 15838 14968 15844 15020
rect 15896 15008 15902 15020
rect 17512 15008 17540 15036
rect 18616 15008 18644 15039
rect 19426 15036 19432 15088
rect 19484 15076 19490 15088
rect 19521 15079 19579 15085
rect 19521 15076 19533 15079
rect 19484 15048 19533 15076
rect 19484 15036 19490 15048
rect 19521 15045 19533 15048
rect 19567 15045 19579 15079
rect 19521 15039 19579 15045
rect 19613 15079 19671 15085
rect 19613 15045 19625 15079
rect 19659 15076 19671 15079
rect 19978 15076 19984 15088
rect 19659 15048 19984 15076
rect 19659 15045 19671 15048
rect 19613 15039 19671 15045
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 15896 14980 18644 15008
rect 19337 15011 19395 15017
rect 15896 14968 15902 14980
rect 19337 14977 19349 15011
rect 19383 15008 19395 15011
rect 19705 15011 19763 15017
rect 19383 14980 19472 15008
rect 19383 14977 19395 14980
rect 19337 14971 19395 14977
rect 19444 14952 19472 14980
rect 19705 14977 19717 15011
rect 19751 15008 19763 15011
rect 20622 15008 20628 15020
rect 19751 14980 20628 15008
rect 19751 14977 19763 14980
rect 19705 14971 19763 14977
rect 16022 14940 16028 14952
rect 15488 14912 16028 14940
rect 16022 14900 16028 14912
rect 16080 14900 16086 14952
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14940 16175 14943
rect 16390 14940 16396 14952
rect 16163 14912 16396 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 16390 14900 16396 14912
rect 16448 14940 16454 14952
rect 17218 14940 17224 14952
rect 16448 14912 17224 14940
rect 16448 14900 16454 14912
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 17494 14900 17500 14952
rect 17552 14900 17558 14952
rect 18598 14900 18604 14952
rect 18656 14940 18662 14952
rect 18693 14943 18751 14949
rect 18693 14940 18705 14943
rect 18656 14912 18705 14940
rect 18656 14900 18662 14912
rect 18693 14909 18705 14912
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 18800 14912 19334 14940
rect 13538 14872 13544 14884
rect 5408 14844 5764 14872
rect 9968 14844 13544 14872
rect 5408 14832 5414 14844
rect 1946 14764 1952 14816
rect 2004 14804 2010 14816
rect 2409 14807 2467 14813
rect 2409 14804 2421 14807
rect 2004 14776 2421 14804
rect 2004 14764 2010 14776
rect 2409 14773 2421 14776
rect 2455 14773 2467 14807
rect 2409 14767 2467 14773
rect 3050 14764 3056 14816
rect 3108 14804 3114 14816
rect 4709 14807 4767 14813
rect 4709 14804 4721 14807
rect 3108 14776 4721 14804
rect 3108 14764 3114 14776
rect 4709 14773 4721 14776
rect 4755 14773 4767 14807
rect 4709 14767 4767 14773
rect 5534 14764 5540 14816
rect 5592 14804 5598 14816
rect 6270 14804 6276 14816
rect 5592 14776 6276 14804
rect 5592 14764 5598 14776
rect 6270 14764 6276 14776
rect 6328 14764 6334 14816
rect 7745 14807 7803 14813
rect 7745 14773 7757 14807
rect 7791 14804 7803 14807
rect 9968 14804 9996 14844
rect 13538 14832 13544 14844
rect 13596 14832 13602 14884
rect 16942 14832 16948 14884
rect 17000 14832 17006 14884
rect 17862 14832 17868 14884
rect 17920 14872 17926 14884
rect 18800 14872 18828 14912
rect 17920 14844 18828 14872
rect 19306 14872 19334 14912
rect 19426 14900 19432 14952
rect 19484 14900 19490 14952
rect 19720 14872 19748 14971
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 22020 15017 22048 15116
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 15008 21235 15011
rect 22005 15011 22063 15017
rect 21223 14980 21680 15008
rect 21223 14977 21235 14980
rect 21177 14971 21235 14977
rect 21358 14900 21364 14952
rect 21416 14900 21422 14952
rect 21652 14940 21680 14980
rect 22005 14977 22017 15011
rect 22051 14977 22063 15011
rect 22112 15008 22140 15116
rect 22922 15104 22928 15156
rect 22980 15144 22986 15156
rect 28821 15147 28879 15153
rect 28821 15144 28833 15147
rect 22980 15116 28833 15144
rect 22980 15104 22986 15116
rect 28821 15113 28833 15116
rect 28867 15113 28879 15147
rect 28821 15107 28879 15113
rect 31205 15147 31263 15153
rect 31205 15113 31217 15147
rect 31251 15144 31263 15147
rect 31662 15144 31668 15156
rect 31251 15116 31668 15144
rect 31251 15113 31263 15116
rect 31205 15107 31263 15113
rect 31662 15104 31668 15116
rect 31720 15104 31726 15156
rect 32674 15144 32680 15156
rect 32232 15116 32680 15144
rect 22186 15036 22192 15088
rect 22244 15076 22250 15088
rect 22244 15048 23152 15076
rect 22244 15036 22250 15048
rect 23124 15017 23152 15048
rect 23290 15036 23296 15088
rect 23348 15076 23354 15088
rect 23385 15079 23443 15085
rect 23385 15076 23397 15079
rect 23348 15048 23397 15076
rect 23348 15036 23354 15048
rect 23385 15045 23397 15048
rect 23431 15045 23443 15079
rect 23385 15039 23443 15045
rect 23934 15036 23940 15088
rect 23992 15036 23998 15088
rect 26234 15036 26240 15088
rect 26292 15076 26298 15088
rect 30837 15079 30895 15085
rect 30837 15076 30849 15079
rect 26292 15048 30849 15076
rect 26292 15036 26298 15048
rect 30837 15045 30849 15048
rect 30883 15045 30895 15079
rect 30837 15039 30895 15045
rect 31053 15079 31111 15085
rect 31053 15045 31065 15079
rect 31099 15076 31111 15079
rect 31386 15076 31392 15088
rect 31099 15048 31392 15076
rect 31099 15045 31111 15048
rect 31053 15039 31111 15045
rect 31386 15036 31392 15048
rect 31444 15036 31450 15088
rect 23109 15011 23167 15017
rect 22112 14980 22324 15008
rect 22005 14971 22063 14977
rect 22094 14940 22100 14952
rect 21652 14912 22100 14940
rect 22094 14900 22100 14912
rect 22152 14900 22158 14952
rect 22189 14943 22247 14949
rect 22189 14909 22201 14943
rect 22235 14909 22247 14943
rect 22296 14940 22324 14980
rect 23109 14977 23121 15011
rect 23155 14977 23167 15011
rect 26786 15008 26792 15020
rect 23109 14971 23167 14977
rect 24596 14980 26792 15008
rect 24596 14940 24624 14980
rect 26786 14968 26792 14980
rect 26844 14968 26850 15020
rect 28258 14968 28264 15020
rect 28316 14968 28322 15020
rect 28442 14968 28448 15020
rect 28500 14968 28506 15020
rect 28534 14968 28540 15020
rect 28592 14968 28598 15020
rect 28634 15011 28692 15017
rect 28634 14977 28646 15011
rect 28680 15008 28692 15011
rect 28810 15008 28816 15020
rect 28680 14980 28816 15008
rect 28680 14977 28692 14980
rect 28634 14971 28692 14977
rect 22296 14912 24624 14940
rect 22189 14903 22247 14909
rect 19306 14844 19748 14872
rect 17920 14832 17926 14844
rect 20622 14832 20628 14884
rect 20680 14872 20686 14884
rect 22204 14872 22232 14903
rect 25130 14900 25136 14952
rect 25188 14900 25194 14952
rect 28350 14900 28356 14952
rect 28408 14940 28414 14952
rect 28644 14940 28672 14971
rect 28810 14968 28816 14980
rect 28868 14968 28874 15020
rect 29086 14968 29092 15020
rect 29144 15008 29150 15020
rect 29365 15011 29423 15017
rect 29365 15008 29377 15011
rect 29144 14980 29377 15008
rect 29144 14968 29150 14980
rect 29365 14977 29377 14980
rect 29411 14977 29423 15011
rect 32232 15008 32260 15116
rect 32674 15104 32680 15116
rect 32732 15104 32738 15156
rect 32858 15104 32864 15156
rect 32916 15144 32922 15156
rect 37829 15147 37887 15153
rect 37829 15144 37841 15147
rect 32916 15116 37841 15144
rect 32916 15104 32922 15116
rect 37829 15113 37841 15116
rect 37875 15113 37887 15147
rect 37829 15107 37887 15113
rect 32582 15036 32588 15088
rect 32640 15076 32646 15088
rect 35066 15076 35072 15088
rect 32640 15048 33074 15076
rect 34900 15048 35072 15076
rect 32640 15036 32646 15048
rect 34900 15020 34928 15048
rect 35066 15036 35072 15048
rect 35124 15036 35130 15088
rect 35158 15036 35164 15088
rect 35216 15036 35222 15088
rect 35894 15036 35900 15088
rect 35952 15036 35958 15088
rect 38470 15036 38476 15088
rect 38528 15036 38534 15088
rect 29365 14971 29423 14977
rect 29932 14980 32260 15008
rect 29932 14952 29960 14980
rect 32306 14968 32312 15020
rect 32364 14968 32370 15020
rect 34882 14968 34888 15020
rect 34940 14968 34946 15020
rect 37737 15011 37795 15017
rect 37737 14977 37749 15011
rect 37783 15008 37795 15011
rect 37826 15008 37832 15020
rect 37783 14980 37832 15008
rect 37783 14977 37795 14980
rect 37737 14971 37795 14977
rect 37826 14968 37832 14980
rect 37884 14968 37890 15020
rect 38654 14968 38660 15020
rect 38712 14968 38718 15020
rect 28408 14912 28672 14940
rect 28408 14900 28414 14912
rect 29914 14900 29920 14952
rect 29972 14900 29978 14952
rect 30282 14900 30288 14952
rect 30340 14940 30346 14952
rect 31018 14940 31024 14952
rect 30340 14912 31024 14940
rect 30340 14900 30346 14912
rect 31018 14900 31024 14912
rect 31076 14940 31082 14952
rect 32324 14940 32352 14968
rect 31076 14912 32352 14940
rect 31076 14900 31082 14912
rect 32582 14900 32588 14952
rect 32640 14900 32646 14952
rect 32674 14900 32680 14952
rect 32732 14940 32738 14952
rect 33962 14940 33968 14952
rect 32732 14912 33968 14940
rect 32732 14900 32738 14912
rect 33962 14900 33968 14912
rect 34020 14900 34026 14952
rect 20680 14844 22232 14872
rect 20680 14832 20686 14844
rect 7791 14776 9996 14804
rect 7791 14773 7803 14776
rect 7745 14767 7803 14773
rect 11238 14764 11244 14816
rect 11296 14804 11302 14816
rect 11606 14804 11612 14816
rect 11296 14776 11612 14804
rect 11296 14764 11302 14776
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 13078 14764 13084 14816
rect 13136 14804 13142 14816
rect 17681 14807 17739 14813
rect 17681 14804 17693 14807
rect 13136 14776 17693 14804
rect 13136 14764 13142 14776
rect 17681 14773 17693 14776
rect 17727 14773 17739 14807
rect 17681 14767 17739 14773
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 19889 14807 19947 14813
rect 19889 14804 19901 14807
rect 18472 14776 19901 14804
rect 18472 14764 18478 14776
rect 19889 14773 19901 14776
rect 19935 14773 19947 14807
rect 19889 14767 19947 14773
rect 20717 14807 20775 14813
rect 20717 14773 20729 14807
rect 20763 14804 20775 14807
rect 21082 14804 21088 14816
rect 20763 14776 21088 14804
rect 20763 14773 20775 14776
rect 20717 14767 20775 14773
rect 21082 14764 21088 14776
rect 21140 14764 21146 14816
rect 26326 14764 26332 14816
rect 26384 14804 26390 14816
rect 28442 14804 28448 14816
rect 26384 14776 28448 14804
rect 26384 14764 26390 14776
rect 28442 14764 28448 14776
rect 28500 14764 28506 14816
rect 31021 14807 31079 14813
rect 31021 14773 31033 14807
rect 31067 14804 31079 14807
rect 31110 14804 31116 14816
rect 31067 14776 31116 14804
rect 31067 14773 31079 14776
rect 31021 14767 31079 14773
rect 31110 14764 31116 14776
rect 31168 14764 31174 14816
rect 31754 14764 31760 14816
rect 31812 14804 31818 14816
rect 34057 14807 34115 14813
rect 34057 14804 34069 14807
rect 31812 14776 34069 14804
rect 31812 14764 31818 14776
rect 34057 14773 34069 14776
rect 34103 14773 34115 14807
rect 34057 14767 34115 14773
rect 36630 14764 36636 14816
rect 36688 14764 36694 14816
rect 1104 14714 39192 14736
rect 1104 14662 5711 14714
rect 5763 14662 5775 14714
rect 5827 14662 5839 14714
rect 5891 14662 5903 14714
rect 5955 14662 5967 14714
rect 6019 14662 15233 14714
rect 15285 14662 15297 14714
rect 15349 14662 15361 14714
rect 15413 14662 15425 14714
rect 15477 14662 15489 14714
rect 15541 14662 24755 14714
rect 24807 14662 24819 14714
rect 24871 14662 24883 14714
rect 24935 14662 24947 14714
rect 24999 14662 25011 14714
rect 25063 14662 34277 14714
rect 34329 14662 34341 14714
rect 34393 14662 34405 14714
rect 34457 14662 34469 14714
rect 34521 14662 34533 14714
rect 34585 14662 39192 14714
rect 1104 14640 39192 14662
rect 1762 14560 1768 14612
rect 1820 14560 1826 14612
rect 2130 14560 2136 14612
rect 2188 14560 2194 14612
rect 2590 14560 2596 14612
rect 2648 14600 2654 14612
rect 2685 14603 2743 14609
rect 2685 14600 2697 14603
rect 2648 14572 2697 14600
rect 2648 14560 2654 14572
rect 2685 14569 2697 14572
rect 2731 14569 2743 14603
rect 2685 14563 2743 14569
rect 4157 14603 4215 14609
rect 4157 14569 4169 14603
rect 4203 14600 4215 14603
rect 4982 14600 4988 14612
rect 4203 14572 4988 14600
rect 4203 14569 4215 14572
rect 4157 14563 4215 14569
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 5092 14572 6684 14600
rect 5092 14532 5120 14572
rect 3344 14504 5120 14532
rect 6656 14532 6684 14572
rect 6730 14560 6736 14612
rect 6788 14600 6794 14612
rect 8754 14600 8760 14612
rect 6788 14572 8760 14600
rect 6788 14560 6794 14572
rect 8754 14560 8760 14572
rect 8812 14560 8818 14612
rect 10321 14603 10379 14609
rect 10321 14569 10333 14603
rect 10367 14600 10379 14603
rect 10367 14572 14320 14600
rect 10367 14569 10379 14572
rect 10321 14563 10379 14569
rect 9214 14532 9220 14544
rect 6656 14504 9220 14532
rect 2314 14424 2320 14476
rect 2372 14464 2378 14476
rect 3050 14464 3056 14476
rect 2372 14436 3056 14464
rect 2372 14424 2378 14436
rect 3050 14424 3056 14436
rect 3108 14464 3114 14476
rect 3344 14473 3372 14504
rect 9214 14492 9220 14504
rect 9272 14492 9278 14544
rect 9950 14532 9956 14544
rect 9508 14504 9956 14532
rect 3145 14467 3203 14473
rect 3145 14464 3157 14467
rect 3108 14436 3157 14464
rect 3108 14424 3114 14436
rect 3145 14433 3157 14436
rect 3191 14433 3203 14467
rect 3145 14427 3203 14433
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4985 14467 5043 14473
rect 4985 14464 4997 14467
rect 4028 14436 4997 14464
rect 4028 14424 4034 14436
rect 4985 14433 4997 14436
rect 5031 14464 5043 14467
rect 7006 14464 7012 14476
rect 5031 14436 7012 14464
rect 5031 14433 5043 14436
rect 4985 14427 5043 14433
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 9508 14464 9536 14504
rect 9950 14492 9956 14504
rect 10008 14492 10014 14544
rect 13262 14532 13268 14544
rect 10796 14504 13268 14532
rect 7116 14436 9536 14464
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14365 1915 14399
rect 1857 14359 1915 14365
rect 1670 14288 1676 14340
rect 1728 14288 1734 14340
rect 1872 14328 1900 14359
rect 1946 14356 1952 14408
rect 2004 14356 2010 14408
rect 3694 14356 3700 14408
rect 3752 14396 3758 14408
rect 4338 14396 4344 14408
rect 3752 14368 4344 14396
rect 3752 14356 3758 14368
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 7116 14396 7144 14436
rect 9582 14424 9588 14476
rect 9640 14424 9646 14476
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14464 9827 14467
rect 10796 14464 10824 14504
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 13446 14492 13452 14544
rect 13504 14532 13510 14544
rect 13725 14535 13783 14541
rect 13725 14532 13737 14535
rect 13504 14504 13737 14532
rect 13504 14492 13510 14504
rect 13725 14501 13737 14504
rect 13771 14501 13783 14535
rect 14292 14532 14320 14572
rect 14550 14560 14556 14612
rect 14608 14600 14614 14612
rect 14608 14572 17448 14600
rect 14608 14560 14614 14572
rect 14292 14504 15056 14532
rect 13725 14495 13783 14501
rect 9815 14436 10824 14464
rect 9815 14433 9827 14436
rect 9769 14427 9827 14433
rect 10870 14424 10876 14476
rect 10928 14424 10934 14476
rect 12710 14464 12716 14476
rect 10980 14436 12716 14464
rect 6394 14368 7144 14396
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 10980 14396 11008 14436
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 15028 14464 15056 14504
rect 16209 14467 16267 14473
rect 16209 14464 16221 14467
rect 13004 14436 13400 14464
rect 15028 14436 16221 14464
rect 7248 14368 11008 14396
rect 7248 14356 7254 14368
rect 11790 14356 11796 14408
rect 11848 14356 11854 14408
rect 11882 14356 11888 14408
rect 11940 14396 11946 14408
rect 13004 14396 13032 14436
rect 11940 14368 13032 14396
rect 11940 14356 11946 14368
rect 13078 14356 13084 14408
rect 13136 14356 13142 14408
rect 13262 14405 13268 14408
rect 13229 14399 13268 14405
rect 13229 14365 13241 14399
rect 13229 14359 13268 14365
rect 13262 14356 13268 14359
rect 13320 14356 13326 14408
rect 13372 14396 13400 14436
rect 16209 14433 16221 14436
rect 16255 14433 16267 14467
rect 16209 14427 16267 14433
rect 13587 14399 13645 14405
rect 13587 14396 13599 14399
rect 13372 14368 13599 14396
rect 13587 14365 13599 14368
rect 13633 14396 13645 14399
rect 13906 14396 13912 14408
rect 13633 14368 13912 14396
rect 13633 14365 13645 14368
rect 13587 14359 13645 14365
rect 13906 14356 13912 14368
rect 13964 14396 13970 14408
rect 14090 14396 14096 14408
rect 13964 14368 14096 14396
rect 13964 14356 13970 14368
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14826 14396 14832 14408
rect 14516 14368 14832 14396
rect 14516 14356 14522 14368
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15930 14396 15936 14408
rect 15068 14368 15936 14396
rect 15068 14356 15074 14368
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 17420 14396 17448 14572
rect 17494 14560 17500 14612
rect 17552 14600 17558 14612
rect 17862 14600 17868 14612
rect 17552 14572 17868 14600
rect 17552 14560 17558 14572
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 19613 14603 19671 14609
rect 19613 14569 19625 14603
rect 19659 14600 19671 14603
rect 19659 14572 26740 14600
rect 19659 14569 19671 14572
rect 19613 14563 19671 14569
rect 18782 14492 18788 14544
rect 18840 14532 18846 14544
rect 18840 14504 20300 14532
rect 18840 14492 18846 14504
rect 17862 14424 17868 14476
rect 17920 14464 17926 14476
rect 20272 14473 20300 14504
rect 22094 14492 22100 14544
rect 22152 14532 22158 14544
rect 22557 14535 22615 14541
rect 22557 14532 22569 14535
rect 22152 14504 22569 14532
rect 22152 14492 22158 14504
rect 22557 14501 22569 14504
rect 22603 14501 22615 14535
rect 26712 14532 26740 14572
rect 26786 14560 26792 14612
rect 26844 14600 26850 14612
rect 38013 14603 38071 14609
rect 38013 14600 38025 14603
rect 26844 14572 38025 14600
rect 26844 14560 26850 14572
rect 38013 14569 38025 14572
rect 38059 14569 38071 14603
rect 38013 14563 38071 14569
rect 27798 14532 27804 14544
rect 26712 14504 27804 14532
rect 22557 14495 22615 14501
rect 27798 14492 27804 14504
rect 27856 14492 27862 14544
rect 27982 14492 27988 14544
rect 28040 14532 28046 14544
rect 28040 14504 29040 14532
rect 28040 14492 28046 14504
rect 29012 14476 29040 14504
rect 32306 14492 32312 14544
rect 32364 14532 32370 14544
rect 34882 14532 34888 14544
rect 32364 14504 34888 14532
rect 32364 14492 32370 14504
rect 34882 14492 34888 14504
rect 34940 14532 34946 14544
rect 34940 14504 35020 14532
rect 34940 14492 34946 14504
rect 20257 14467 20315 14473
rect 17920 14436 19334 14464
rect 17920 14424 17926 14436
rect 18417 14399 18475 14405
rect 18417 14396 18429 14399
rect 17420 14368 18429 14396
rect 18417 14365 18429 14368
rect 18463 14365 18475 14399
rect 18417 14359 18475 14365
rect 3053 14331 3111 14337
rect 1872 14300 2774 14328
rect 2746 14260 2774 14300
rect 3053 14297 3065 14331
rect 3099 14328 3111 14331
rect 3142 14328 3148 14340
rect 3099 14300 3148 14328
rect 3099 14297 3111 14300
rect 3053 14291 3111 14297
rect 3142 14288 3148 14300
rect 3200 14288 3206 14340
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 3973 14331 4031 14337
rect 3973 14328 3985 14331
rect 3660 14300 3985 14328
rect 3660 14288 3666 14300
rect 3973 14297 3985 14300
rect 4019 14297 4031 14331
rect 3973 14291 4031 14297
rect 4189 14331 4247 14337
rect 4189 14297 4201 14331
rect 4235 14328 4247 14331
rect 5166 14328 5172 14340
rect 4235 14300 5172 14328
rect 4235 14297 4247 14300
rect 4189 14291 4247 14297
rect 5166 14288 5172 14300
rect 5224 14288 5230 14340
rect 5261 14331 5319 14337
rect 5261 14297 5273 14331
rect 5307 14297 5319 14331
rect 5261 14291 5319 14297
rect 4341 14263 4399 14269
rect 4341 14260 4353 14263
rect 2746 14232 4353 14260
rect 4341 14229 4353 14232
rect 4387 14229 4399 14263
rect 5283 14260 5311 14291
rect 6546 14288 6552 14340
rect 6604 14328 6610 14340
rect 7929 14331 7987 14337
rect 7929 14328 7941 14331
rect 6604 14300 7941 14328
rect 6604 14288 6610 14300
rect 7929 14297 7941 14300
rect 7975 14297 7987 14331
rect 8938 14328 8944 14340
rect 7929 14291 7987 14297
rect 8036 14300 8944 14328
rect 6638 14260 6644 14272
rect 5283 14232 6644 14260
rect 4341 14223 4399 14229
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 6730 14220 6736 14272
rect 6788 14220 6794 14272
rect 7098 14220 7104 14272
rect 7156 14260 7162 14272
rect 8036 14260 8064 14300
rect 8938 14288 8944 14300
rect 8996 14288 9002 14340
rect 10689 14331 10747 14337
rect 10689 14297 10701 14331
rect 10735 14328 10747 14331
rect 12066 14328 12072 14340
rect 10735 14300 12072 14328
rect 10735 14297 10747 14300
rect 10689 14291 10747 14297
rect 12066 14288 12072 14300
rect 12124 14288 12130 14340
rect 12250 14288 12256 14340
rect 12308 14288 12314 14340
rect 12986 14288 12992 14340
rect 13044 14328 13050 14340
rect 13357 14331 13415 14337
rect 13357 14328 13369 14331
rect 13044 14300 13369 14328
rect 13044 14288 13050 14300
rect 13357 14297 13369 14300
rect 13403 14297 13415 14331
rect 13357 14291 13415 14297
rect 13446 14288 13452 14340
rect 13504 14288 13510 14340
rect 15381 14331 15439 14337
rect 15381 14297 15393 14331
rect 15427 14328 15439 14331
rect 15654 14328 15660 14340
rect 15427 14300 15660 14328
rect 15427 14297 15439 14300
rect 15381 14291 15439 14297
rect 15654 14288 15660 14300
rect 15712 14328 15718 14340
rect 16206 14328 16212 14340
rect 15712 14300 16212 14328
rect 15712 14288 15718 14300
rect 16206 14288 16212 14300
rect 16264 14288 16270 14340
rect 16666 14288 16672 14340
rect 16724 14288 16730 14340
rect 17586 14328 17592 14340
rect 17512 14300 17592 14328
rect 7156 14232 8064 14260
rect 7156 14220 7162 14232
rect 8570 14220 8576 14272
rect 8628 14260 8634 14272
rect 9125 14263 9183 14269
rect 9125 14260 9137 14263
rect 8628 14232 9137 14260
rect 8628 14220 8634 14232
rect 9125 14229 9137 14232
rect 9171 14229 9183 14263
rect 9125 14223 9183 14229
rect 9490 14220 9496 14272
rect 9548 14220 9554 14272
rect 10781 14263 10839 14269
rect 10781 14229 10793 14263
rect 10827 14260 10839 14263
rect 17512 14260 17540 14300
rect 17586 14288 17592 14300
rect 17644 14328 17650 14340
rect 17957 14331 18015 14337
rect 17957 14328 17969 14331
rect 17644 14300 17969 14328
rect 17644 14288 17650 14300
rect 17957 14297 17969 14300
rect 18003 14297 18015 14331
rect 17957 14291 18015 14297
rect 18506 14288 18512 14340
rect 18564 14328 18570 14340
rect 18693 14331 18751 14337
rect 18693 14328 18705 14331
rect 18564 14300 18705 14328
rect 18564 14288 18570 14300
rect 18693 14297 18705 14300
rect 18739 14297 18751 14331
rect 18693 14291 18751 14297
rect 10827 14232 17540 14260
rect 19306 14260 19334 14436
rect 20257 14433 20269 14467
rect 20303 14464 20315 14467
rect 20622 14464 20628 14476
rect 20303 14436 20628 14464
rect 20303 14433 20315 14436
rect 20257 14427 20315 14433
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 25041 14467 25099 14473
rect 25041 14464 25053 14467
rect 24912 14436 25053 14464
rect 24912 14424 24918 14436
rect 25041 14433 25053 14436
rect 25087 14464 25099 14467
rect 25314 14464 25320 14476
rect 25087 14436 25320 14464
rect 25087 14433 25099 14436
rect 25041 14427 25099 14433
rect 25314 14424 25320 14436
rect 25372 14424 25378 14476
rect 27614 14424 27620 14476
rect 27672 14464 27678 14476
rect 28902 14464 28908 14476
rect 27672 14436 28908 14464
rect 27672 14424 27678 14436
rect 28902 14424 28908 14436
rect 28960 14424 28966 14476
rect 28994 14424 29000 14476
rect 29052 14424 29058 14476
rect 29270 14424 29276 14476
rect 29328 14464 29334 14476
rect 30285 14467 30343 14473
rect 30285 14464 30297 14467
rect 29328 14436 30297 14464
rect 29328 14424 29334 14436
rect 30285 14433 30297 14436
rect 30331 14464 30343 14467
rect 30466 14464 30472 14476
rect 30331 14436 30472 14464
rect 30331 14433 30343 14436
rect 30285 14427 30343 14433
rect 30466 14424 30472 14436
rect 30524 14424 30530 14476
rect 31018 14424 31024 14476
rect 31076 14424 31082 14476
rect 34992 14473 35020 14504
rect 37366 14492 37372 14544
rect 37424 14492 37430 14544
rect 34977 14467 35035 14473
rect 34977 14433 34989 14467
rect 35023 14433 35035 14467
rect 34977 14427 35035 14433
rect 19886 14356 19892 14408
rect 19944 14396 19950 14408
rect 19981 14399 20039 14405
rect 19981 14396 19993 14399
rect 19944 14368 19993 14396
rect 19944 14356 19950 14368
rect 19981 14365 19993 14368
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 20809 14399 20867 14405
rect 20809 14396 20821 14399
rect 20772 14368 20821 14396
rect 20772 14356 20778 14368
rect 20809 14365 20821 14368
rect 20855 14365 20867 14399
rect 20809 14359 20867 14365
rect 27801 14399 27859 14405
rect 27801 14365 27813 14399
rect 27847 14396 27859 14399
rect 30190 14396 30196 14408
rect 27847 14368 30196 14396
rect 27847 14365 27859 14368
rect 27801 14359 27859 14365
rect 30190 14356 30196 14368
rect 30248 14356 30254 14408
rect 33134 14356 33140 14408
rect 33192 14396 33198 14408
rect 33413 14399 33471 14405
rect 33413 14396 33425 14399
rect 33192 14368 33425 14396
rect 33192 14356 33198 14368
rect 33413 14365 33425 14368
rect 33459 14365 33471 14399
rect 33413 14359 33471 14365
rect 33502 14356 33508 14408
rect 33560 14396 33566 14408
rect 33781 14399 33839 14405
rect 33781 14396 33793 14399
rect 33560 14368 33793 14396
rect 33560 14356 33566 14368
rect 33781 14365 33793 14368
rect 33827 14365 33839 14399
rect 33781 14359 33839 14365
rect 36354 14356 36360 14408
rect 36412 14356 36418 14408
rect 37182 14356 37188 14408
rect 37240 14356 37246 14408
rect 37921 14399 37979 14405
rect 37921 14365 37933 14399
rect 37967 14396 37979 14399
rect 38102 14396 38108 14408
rect 37967 14368 38108 14396
rect 37967 14365 37979 14368
rect 37921 14359 37979 14365
rect 38102 14356 38108 14368
rect 38160 14356 38166 14408
rect 21082 14288 21088 14340
rect 21140 14288 21146 14340
rect 21174 14288 21180 14340
rect 21232 14328 21238 14340
rect 21232 14300 21574 14328
rect 21232 14288 21238 14300
rect 23658 14288 23664 14340
rect 23716 14328 23722 14340
rect 25317 14331 25375 14337
rect 25317 14328 25329 14331
rect 23716 14300 25329 14328
rect 23716 14288 23722 14300
rect 25317 14297 25329 14300
rect 25363 14297 25375 14331
rect 27893 14331 27951 14337
rect 26542 14300 26648 14328
rect 25317 14291 25375 14297
rect 20073 14263 20131 14269
rect 20073 14260 20085 14263
rect 19306 14232 20085 14260
rect 10827 14229 10839 14232
rect 10781 14223 10839 14229
rect 20073 14229 20085 14232
rect 20119 14260 20131 14263
rect 23842 14260 23848 14272
rect 20119 14232 23848 14260
rect 20119 14229 20131 14232
rect 20073 14223 20131 14229
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 26620 14260 26648 14300
rect 27893 14297 27905 14331
rect 27939 14328 27951 14331
rect 28718 14328 28724 14340
rect 27939 14300 28724 14328
rect 27939 14297 27951 14300
rect 27893 14291 27951 14297
rect 28718 14288 28724 14300
rect 28776 14288 28782 14340
rect 28813 14331 28871 14337
rect 28813 14297 28825 14331
rect 28859 14328 28871 14331
rect 29914 14328 29920 14340
rect 28859 14300 29920 14328
rect 28859 14297 28871 14300
rect 28813 14291 28871 14297
rect 29914 14288 29920 14300
rect 29972 14288 29978 14340
rect 30101 14331 30159 14337
rect 30101 14297 30113 14331
rect 30147 14328 30159 14331
rect 30742 14328 30748 14340
rect 30147 14300 30748 14328
rect 30147 14297 30159 14300
rect 30101 14291 30159 14297
rect 30742 14288 30748 14300
rect 30800 14288 30806 14340
rect 31294 14288 31300 14340
rect 31352 14288 31358 14340
rect 32522 14300 33916 14328
rect 26694 14260 26700 14272
rect 26620 14232 26700 14260
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 26786 14220 26792 14272
rect 26844 14220 26850 14272
rect 28442 14220 28448 14272
rect 28500 14220 28506 14272
rect 28994 14220 29000 14272
rect 29052 14260 29058 14272
rect 29270 14260 29276 14272
rect 29052 14232 29276 14260
rect 29052 14220 29058 14232
rect 29270 14220 29276 14232
rect 29328 14220 29334 14272
rect 29733 14263 29791 14269
rect 29733 14229 29745 14263
rect 29779 14260 29791 14263
rect 30006 14260 30012 14272
rect 29779 14232 30012 14260
rect 29779 14229 29791 14232
rect 29733 14223 29791 14229
rect 30006 14220 30012 14232
rect 30064 14220 30070 14272
rect 30193 14263 30251 14269
rect 30193 14229 30205 14263
rect 30239 14260 30251 14263
rect 31478 14260 31484 14272
rect 30239 14232 31484 14260
rect 30239 14229 30251 14232
rect 30193 14223 30251 14229
rect 31478 14220 31484 14232
rect 31536 14220 31542 14272
rect 31570 14220 31576 14272
rect 31628 14260 31634 14272
rect 32769 14263 32827 14269
rect 32769 14260 32781 14263
rect 31628 14232 32781 14260
rect 31628 14220 31634 14232
rect 32769 14229 32781 14232
rect 32815 14229 32827 14263
rect 33888 14260 33916 14300
rect 35250 14288 35256 14340
rect 35308 14288 35314 14340
rect 36630 14260 36636 14272
rect 33888 14232 36636 14260
rect 32769 14223 32827 14229
rect 36630 14220 36636 14232
rect 36688 14220 36694 14272
rect 36722 14220 36728 14272
rect 36780 14220 36786 14272
rect 1104 14170 39352 14192
rect 1104 14118 10472 14170
rect 10524 14118 10536 14170
rect 10588 14118 10600 14170
rect 10652 14118 10664 14170
rect 10716 14118 10728 14170
rect 10780 14118 19994 14170
rect 20046 14118 20058 14170
rect 20110 14118 20122 14170
rect 20174 14118 20186 14170
rect 20238 14118 20250 14170
rect 20302 14118 29516 14170
rect 29568 14118 29580 14170
rect 29632 14118 29644 14170
rect 29696 14118 29708 14170
rect 29760 14118 29772 14170
rect 29824 14118 39038 14170
rect 39090 14118 39102 14170
rect 39154 14118 39166 14170
rect 39218 14118 39230 14170
rect 39282 14118 39294 14170
rect 39346 14118 39352 14170
rect 1104 14096 39352 14118
rect 6546 14056 6552 14068
rect 4172 14028 6552 14056
rect 2038 13948 2044 14000
rect 2096 13948 2102 14000
rect 3418 13988 3424 14000
rect 3266 13960 3424 13988
rect 3418 13948 3424 13960
rect 3476 13948 3482 14000
rect 4172 13988 4200 14028
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 8297 14059 8355 14065
rect 8297 14056 8309 14059
rect 6696 14028 8309 14056
rect 6696 14016 6702 14028
rect 8297 14025 8309 14028
rect 8343 14025 8355 14059
rect 8297 14019 8355 14025
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8665 14059 8723 14065
rect 8665 14056 8677 14059
rect 8536 14028 8677 14056
rect 8536 14016 8542 14028
rect 8665 14025 8677 14028
rect 8711 14025 8723 14059
rect 8665 14019 8723 14025
rect 10781 14059 10839 14065
rect 10781 14025 10793 14059
rect 10827 14056 10839 14059
rect 11606 14056 11612 14068
rect 10827 14028 11612 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 14550 14056 14556 14068
rect 12836 14028 14556 14056
rect 4080 13960 4200 13988
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 4080 13929 4108 13960
rect 10042 13948 10048 14000
rect 10100 13988 10106 14000
rect 10413 13991 10471 13997
rect 10413 13988 10425 13991
rect 10100 13960 10425 13988
rect 10100 13948 10106 13960
rect 10413 13957 10425 13960
rect 10459 13957 10471 13991
rect 10413 13951 10471 13957
rect 10629 13991 10687 13997
rect 10629 13957 10641 13991
rect 10675 13988 10687 13991
rect 12836 13988 12864 14028
rect 14550 14016 14556 14028
rect 14608 14016 14614 14068
rect 15010 14056 15016 14068
rect 14660 14028 15016 14056
rect 14366 13988 14372 14000
rect 10675 13960 12864 13988
rect 14214 13960 14372 13988
rect 10675 13957 10687 13960
rect 10629 13951 10687 13957
rect 14366 13948 14372 13960
rect 14424 13948 14430 14000
rect 14458 13948 14464 14000
rect 14516 13988 14522 14000
rect 14660 13988 14688 14028
rect 15010 14016 15016 14028
rect 15068 14056 15074 14068
rect 25222 14056 25228 14068
rect 15068 14028 25228 14056
rect 15068 14016 15074 14028
rect 14516 13960 14688 13988
rect 14516 13948 14522 13960
rect 15102 13948 15108 14000
rect 15160 13988 15166 14000
rect 15562 13988 15568 14000
rect 15160 13960 15568 13988
rect 15160 13948 15166 13960
rect 15562 13948 15568 13960
rect 15620 13948 15626 14000
rect 16209 13991 16267 13997
rect 16209 13957 16221 13991
rect 16255 13988 16267 13991
rect 16666 13988 16672 14000
rect 16255 13960 16672 13988
rect 16255 13957 16267 13960
rect 16209 13951 16267 13957
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 17586 13948 17592 14000
rect 17644 13988 17650 14000
rect 17644 13960 19334 13988
rect 17644 13948 17650 13960
rect 4065 13923 4123 13929
rect 4065 13920 4077 13923
rect 4028 13892 4077 13920
rect 4028 13880 4034 13892
rect 4065 13889 4077 13892
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 5442 13880 5448 13932
rect 5500 13880 5506 13932
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 1765 13855 1823 13861
rect 1765 13821 1777 13855
rect 1811 13852 1823 13855
rect 2130 13852 2136 13864
rect 1811 13824 2136 13852
rect 1811 13821 1823 13824
rect 1765 13815 1823 13821
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 3513 13855 3571 13861
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 3694 13852 3700 13864
rect 3559 13824 3700 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3694 13812 3700 13824
rect 3752 13812 3758 13864
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 5813 13855 5871 13861
rect 5813 13852 5825 13855
rect 5592 13824 5825 13852
rect 5592 13812 5598 13824
rect 5813 13821 5825 13824
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 4062 13676 4068 13728
rect 4120 13716 4126 13728
rect 4322 13719 4380 13725
rect 4322 13716 4334 13719
rect 4120 13688 4334 13716
rect 4120 13676 4126 13688
rect 4322 13685 4334 13688
rect 4368 13685 4380 13719
rect 4322 13679 4380 13685
rect 5626 13676 5632 13728
rect 5684 13716 5690 13728
rect 6638 13716 6644 13728
rect 5684 13688 6644 13716
rect 5684 13676 5690 13688
rect 6638 13676 6644 13688
rect 6696 13676 6702 13728
rect 6932 13716 6960 13883
rect 8018 13880 8024 13932
rect 8076 13920 8082 13932
rect 8757 13923 8815 13929
rect 8757 13920 8769 13923
rect 8076 13892 8769 13920
rect 8076 13880 8082 13892
rect 8757 13889 8769 13892
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 8996 13892 9505 13920
rect 8996 13880 9002 13892
rect 9493 13889 9505 13892
rect 9539 13920 9551 13923
rect 10502 13920 10508 13932
rect 9539 13892 10508 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 11974 13880 11980 13932
rect 12032 13880 12038 13932
rect 12618 13880 12624 13932
rect 12676 13920 12682 13932
rect 12713 13923 12771 13929
rect 12713 13920 12725 13923
rect 12676 13892 12725 13920
rect 12676 13880 12682 13892
rect 12713 13889 12725 13892
rect 12759 13889 12771 13923
rect 14642 13920 14648 13932
rect 12713 13883 12771 13889
rect 14200 13892 14648 13920
rect 7006 13812 7012 13864
rect 7064 13852 7070 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7064 13824 7757 13852
rect 7064 13812 7070 13824
rect 7745 13821 7757 13824
rect 7791 13852 7803 13855
rect 8294 13852 8300 13864
rect 7791 13824 8300 13852
rect 7791 13821 7803 13824
rect 7745 13815 7803 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 9815 13824 9849 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 8202 13744 8208 13796
rect 8260 13784 8266 13796
rect 8864 13784 8892 13815
rect 9784 13784 9812 13815
rect 13446 13812 13452 13864
rect 13504 13852 13510 13864
rect 14200 13852 14228 13892
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13889 15347 13923
rect 15289 13883 15347 13889
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 16117 13923 16175 13929
rect 15427 13892 15792 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 13504 13824 14228 13852
rect 14461 13855 14519 13861
rect 13504 13812 13510 13824
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 14826 13852 14832 13864
rect 14507 13824 14832 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 14826 13812 14832 13824
rect 14884 13852 14890 13864
rect 15304 13852 15332 13883
rect 14884 13824 15332 13852
rect 14884 13812 14890 13824
rect 15562 13812 15568 13864
rect 15620 13812 15626 13864
rect 10318 13784 10324 13796
rect 8260 13756 8892 13784
rect 9600 13756 10324 13784
rect 8260 13744 8266 13756
rect 7190 13716 7196 13728
rect 6932 13688 7196 13716
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 8018 13676 8024 13728
rect 8076 13716 8082 13728
rect 9600 13716 9628 13756
rect 10318 13744 10324 13756
rect 10376 13744 10382 13796
rect 10502 13744 10508 13796
rect 10560 13784 10566 13796
rect 12526 13784 12532 13796
rect 10560 13756 12532 13784
rect 10560 13744 10566 13756
rect 10612 13725 10640 13756
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 14921 13787 14979 13793
rect 14921 13784 14933 13787
rect 14016 13756 14933 13784
rect 8076 13688 9628 13716
rect 10597 13719 10655 13725
rect 8076 13676 8082 13688
rect 10597 13685 10609 13719
rect 10643 13685 10655 13719
rect 10597 13679 10655 13685
rect 12066 13676 12072 13728
rect 12124 13676 12130 13728
rect 12976 13719 13034 13725
rect 12976 13685 12988 13719
rect 13022 13716 13034 13719
rect 14016 13716 14044 13756
rect 14921 13753 14933 13756
rect 14967 13753 14979 13787
rect 14921 13747 14979 13753
rect 13022 13688 14044 13716
rect 13022 13685 13034 13688
rect 12976 13679 13034 13685
rect 14642 13676 14648 13728
rect 14700 13716 14706 13728
rect 15102 13716 15108 13728
rect 14700 13688 15108 13716
rect 14700 13676 14706 13688
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 15764 13716 15792 13892
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16390 13920 16396 13932
rect 16163 13892 16396 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 17221 13923 17279 13929
rect 17221 13889 17233 13923
rect 17267 13920 17279 13923
rect 18230 13920 18236 13932
rect 17267 13892 18236 13920
rect 17267 13889 17279 13892
rect 17221 13883 17279 13889
rect 16666 13812 16672 13864
rect 16724 13852 16730 13864
rect 17236 13852 17264 13883
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 19306 13920 19334 13960
rect 19702 13948 19708 14000
rect 19760 13948 19766 14000
rect 20714 13948 20720 14000
rect 20772 13988 20778 14000
rect 21082 13988 21088 14000
rect 20772 13960 21088 13988
rect 20772 13948 20778 13960
rect 21082 13948 21088 13960
rect 21140 13948 21146 14000
rect 21468 13997 21496 14028
rect 25222 14016 25228 14028
rect 25280 14016 25286 14068
rect 27890 14056 27896 14068
rect 25332 14028 27896 14056
rect 21453 13991 21511 13997
rect 21453 13957 21465 13991
rect 21499 13957 21511 13991
rect 21453 13951 21511 13957
rect 23474 13948 23480 14000
rect 23532 13948 23538 14000
rect 23842 13948 23848 14000
rect 23900 13988 23906 14000
rect 25332 13988 25360 14028
rect 27890 14016 27896 14028
rect 27948 14016 27954 14068
rect 29362 14056 29368 14068
rect 28184 14028 29368 14056
rect 23900 13960 25360 13988
rect 26358 13960 28120 13988
rect 23900 13948 23906 13960
rect 20438 13920 20444 13932
rect 19306 13892 20444 13920
rect 18601 13883 18659 13889
rect 16724 13824 17264 13852
rect 17313 13855 17371 13861
rect 16724 13812 16730 13824
rect 17313 13821 17325 13855
rect 17359 13821 17371 13855
rect 17313 13815 17371 13821
rect 17218 13744 17224 13796
rect 17276 13784 17282 13796
rect 17328 13784 17356 13815
rect 17402 13812 17408 13864
rect 17460 13812 17466 13864
rect 17276 13756 17356 13784
rect 17420 13784 17448 13812
rect 18230 13784 18236 13796
rect 17420 13756 18236 13784
rect 17276 13744 17282 13756
rect 16666 13716 16672 13728
rect 15712 13688 16672 13716
rect 15712 13676 15718 13688
rect 16666 13676 16672 13688
rect 16724 13676 16730 13728
rect 16850 13676 16856 13728
rect 16908 13676 16914 13728
rect 17328 13716 17356 13756
rect 18230 13744 18236 13756
rect 18288 13784 18294 13796
rect 18616 13784 18644 13883
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 20732 13892 21312 13920
rect 19153 13855 19211 13861
rect 19153 13821 19165 13855
rect 19199 13852 19211 13855
rect 20622 13852 20628 13864
rect 19199 13824 20628 13852
rect 19199 13821 19211 13824
rect 19153 13815 19211 13821
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 18782 13784 18788 13796
rect 18288 13756 18788 13784
rect 18288 13744 18294 13756
rect 18782 13744 18788 13756
rect 18840 13744 18846 13796
rect 19426 13744 19432 13796
rect 19484 13784 19490 13796
rect 20732 13784 20760 13892
rect 21284 13852 21312 13892
rect 21358 13880 21364 13932
rect 21416 13920 21422 13932
rect 21634 13920 21640 13932
rect 21416 13892 21640 13920
rect 21416 13880 21422 13892
rect 21634 13880 21640 13892
rect 21692 13880 21698 13932
rect 22186 13880 22192 13932
rect 22244 13880 22250 13932
rect 24854 13880 24860 13932
rect 24912 13880 24918 13932
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13920 27215 13923
rect 27430 13920 27436 13932
rect 27203 13892 27436 13920
rect 27203 13889 27215 13892
rect 27157 13883 27215 13889
rect 27430 13880 27436 13892
rect 27488 13880 27494 13932
rect 23937 13855 23995 13861
rect 23937 13852 23949 13855
rect 19484 13756 20760 13784
rect 21008 13824 21220 13852
rect 21284 13824 23949 13852
rect 19484 13744 19490 13756
rect 17678 13716 17684 13728
rect 17328 13688 17684 13716
rect 17678 13676 17684 13688
rect 17736 13676 17742 13728
rect 17770 13676 17776 13728
rect 17828 13716 17834 13728
rect 21008 13716 21036 13824
rect 21192 13784 21220 13824
rect 23937 13821 23949 13824
rect 23983 13821 23995 13855
rect 24872 13852 24900 13880
rect 25130 13852 25136 13864
rect 24872 13824 25136 13852
rect 23937 13815 23995 13821
rect 25130 13812 25136 13824
rect 25188 13812 25194 13864
rect 27246 13812 27252 13864
rect 27304 13812 27310 13864
rect 28092 13852 28120 13960
rect 28184 13929 28212 14028
rect 29362 14016 29368 14028
rect 29420 14016 29426 14068
rect 29914 14016 29920 14068
rect 29972 14056 29978 14068
rect 30374 14056 30380 14068
rect 29972 14028 30380 14056
rect 29972 14016 29978 14028
rect 30374 14016 30380 14028
rect 30432 14016 30438 14068
rect 30834 14016 30840 14068
rect 30892 14056 30898 14068
rect 32309 14059 32367 14065
rect 32309 14056 32321 14059
rect 30892 14028 32321 14056
rect 30892 14016 30898 14028
rect 32309 14025 32321 14028
rect 32355 14025 32367 14059
rect 32309 14019 32367 14025
rect 32674 14016 32680 14068
rect 32732 14056 32738 14068
rect 33686 14056 33692 14068
rect 32732 14028 33692 14056
rect 32732 14016 32738 14028
rect 33686 14016 33692 14028
rect 33744 14016 33750 14068
rect 34149 14059 34207 14065
rect 34149 14025 34161 14059
rect 34195 14056 34207 14059
rect 34606 14056 34612 14068
rect 34195 14028 34612 14056
rect 34195 14025 34207 14028
rect 34149 14019 34207 14025
rect 34606 14016 34612 14028
rect 34664 14016 34670 14068
rect 34698 14016 34704 14068
rect 34756 14016 34762 14068
rect 35250 14016 35256 14068
rect 35308 14056 35314 14068
rect 35437 14059 35495 14065
rect 35437 14056 35449 14059
rect 35308 14028 35449 14056
rect 35308 14016 35314 14028
rect 35437 14025 35449 14028
rect 35483 14025 35495 14059
rect 35437 14019 35495 14025
rect 35805 14059 35863 14065
rect 35805 14025 35817 14059
rect 35851 14056 35863 14059
rect 36722 14056 36728 14068
rect 35851 14028 36728 14056
rect 35851 14025 35863 14028
rect 35805 14019 35863 14025
rect 28442 13948 28448 14000
rect 28500 13948 28506 14000
rect 28718 13948 28724 14000
rect 28776 13988 28782 14000
rect 33318 13988 33324 14000
rect 28776 13960 28934 13988
rect 31312 13960 33324 13988
rect 28776 13948 28782 13960
rect 28169 13923 28227 13929
rect 28169 13889 28181 13923
rect 28215 13889 28227 13923
rect 28169 13883 28227 13889
rect 30190 13880 30196 13932
rect 30248 13920 30254 13932
rect 31312 13929 31340 13960
rect 33318 13948 33324 13960
rect 33376 13948 33382 14000
rect 33704 13988 33732 14016
rect 33781 13991 33839 13997
rect 33781 13988 33793 13991
rect 33704 13960 33793 13988
rect 33781 13957 33793 13960
rect 33827 13957 33839 13991
rect 33781 13951 33839 13957
rect 34238 13948 34244 14000
rect 34296 13988 34302 14000
rect 35820 13988 35848 14019
rect 36722 14016 36728 14028
rect 36780 14016 36786 14068
rect 34296 13960 35848 13988
rect 34296 13948 34302 13960
rect 36630 13948 36636 14000
rect 36688 13988 36694 14000
rect 37553 13991 37611 13997
rect 37553 13988 37565 13991
rect 36688 13960 37565 13988
rect 36688 13948 36694 13960
rect 37553 13957 37565 13960
rect 37599 13957 37611 13991
rect 37553 13951 37611 13957
rect 30561 13923 30619 13929
rect 30561 13920 30573 13923
rect 30248 13892 30573 13920
rect 30248 13880 30254 13892
rect 30561 13889 30573 13892
rect 30607 13889 30619 13923
rect 30561 13883 30619 13889
rect 31297 13923 31355 13929
rect 31297 13889 31309 13923
rect 31343 13889 31355 13923
rect 31297 13883 31355 13889
rect 32677 13923 32735 13929
rect 32677 13889 32689 13923
rect 32723 13920 32735 13923
rect 33042 13920 33048 13932
rect 32723 13892 33048 13920
rect 32723 13889 32735 13892
rect 32677 13883 32735 13889
rect 33042 13880 33048 13892
rect 33100 13880 33106 13932
rect 33597 13923 33655 13929
rect 33597 13889 33609 13923
rect 33643 13920 33655 13923
rect 33686 13920 33692 13932
rect 33643 13892 33692 13920
rect 33643 13889 33655 13892
rect 33597 13883 33655 13889
rect 33686 13880 33692 13892
rect 33744 13880 33750 13932
rect 33873 13923 33931 13929
rect 33873 13889 33885 13923
rect 33919 13889 33931 13923
rect 33873 13883 33931 13889
rect 30653 13855 30711 13861
rect 30653 13852 30665 13855
rect 28092 13824 30665 13852
rect 30653 13821 30665 13824
rect 30699 13821 30711 13855
rect 31846 13852 31852 13864
rect 30653 13815 30711 13821
rect 31404 13824 31852 13852
rect 21818 13784 21824 13796
rect 21192 13756 21824 13784
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 17828 13688 21036 13716
rect 17828 13676 17834 13688
rect 21082 13676 21088 13728
rect 21140 13716 21146 13728
rect 22186 13716 22192 13728
rect 21140 13688 22192 13716
rect 21140 13676 21146 13688
rect 22186 13676 22192 13688
rect 22244 13676 22250 13728
rect 22462 13725 22468 13728
rect 22452 13719 22468 13725
rect 22452 13685 22464 13719
rect 22452 13679 22468 13685
rect 22462 13676 22468 13679
rect 22520 13676 22526 13728
rect 25120 13719 25178 13725
rect 25120 13685 25132 13719
rect 25166 13716 25178 13719
rect 25866 13716 25872 13728
rect 25166 13688 25872 13716
rect 25166 13685 25178 13688
rect 25120 13679 25178 13685
rect 25866 13676 25872 13688
rect 25924 13676 25930 13728
rect 26510 13676 26516 13728
rect 26568 13716 26574 13728
rect 26605 13719 26663 13725
rect 26605 13716 26617 13719
rect 26568 13688 26617 13716
rect 26568 13676 26574 13688
rect 26605 13685 26617 13688
rect 26651 13685 26663 13719
rect 26605 13679 26663 13685
rect 28074 13676 28080 13728
rect 28132 13716 28138 13728
rect 28902 13716 28908 13728
rect 28132 13688 28908 13716
rect 28132 13676 28138 13688
rect 28902 13676 28908 13688
rect 28960 13676 28966 13728
rect 31404 13725 31432 13824
rect 31846 13812 31852 13824
rect 31904 13812 31910 13864
rect 32766 13812 32772 13864
rect 32824 13812 32830 13864
rect 32953 13855 33011 13861
rect 32953 13821 32965 13855
rect 32999 13852 33011 13855
rect 33134 13852 33140 13864
rect 32999 13824 33140 13852
rect 32999 13821 33011 13824
rect 32953 13815 33011 13821
rect 33134 13812 33140 13824
rect 33192 13852 33198 13864
rect 33502 13852 33508 13864
rect 33192 13824 33508 13852
rect 33192 13812 33198 13824
rect 33502 13812 33508 13824
rect 33560 13812 33566 13864
rect 33888 13784 33916 13883
rect 33962 13880 33968 13932
rect 34020 13880 34026 13932
rect 34609 13923 34667 13929
rect 34609 13889 34621 13923
rect 34655 13920 34667 13923
rect 35066 13920 35072 13932
rect 34655 13892 35072 13920
rect 34655 13889 34667 13892
rect 34609 13883 34667 13889
rect 35066 13880 35072 13892
rect 35124 13880 35130 13932
rect 36725 13923 36783 13929
rect 36725 13889 36737 13923
rect 36771 13920 36783 13923
rect 37461 13923 37519 13929
rect 36771 13892 37412 13920
rect 36771 13889 36783 13892
rect 36725 13883 36783 13889
rect 35894 13812 35900 13864
rect 35952 13812 35958 13864
rect 35989 13855 36047 13861
rect 35989 13821 36001 13855
rect 36035 13821 36047 13855
rect 35989 13815 36047 13821
rect 34238 13784 34244 13796
rect 33888 13756 34244 13784
rect 34238 13744 34244 13756
rect 34296 13744 34302 13796
rect 35710 13744 35716 13796
rect 35768 13784 35774 13796
rect 36004 13784 36032 13815
rect 36814 13812 36820 13864
rect 36872 13812 36878 13864
rect 37384 13852 37412 13892
rect 37461 13889 37473 13923
rect 37507 13920 37519 13923
rect 38102 13920 38108 13932
rect 37507 13892 38108 13920
rect 37507 13889 37519 13892
rect 37461 13883 37519 13889
rect 38102 13880 38108 13892
rect 38160 13880 38166 13932
rect 37826 13852 37832 13864
rect 37384 13824 37832 13852
rect 37826 13812 37832 13824
rect 37884 13812 37890 13864
rect 35768 13756 36032 13784
rect 35768 13744 35774 13756
rect 36446 13744 36452 13796
rect 36504 13784 36510 13796
rect 37274 13784 37280 13796
rect 36504 13756 37280 13784
rect 36504 13744 36510 13756
rect 37274 13744 37280 13756
rect 37332 13744 37338 13796
rect 31389 13719 31447 13725
rect 31389 13685 31401 13719
rect 31435 13685 31447 13719
rect 31389 13679 31447 13685
rect 33042 13676 33048 13728
rect 33100 13716 33106 13728
rect 35618 13716 35624 13728
rect 33100 13688 35624 13716
rect 33100 13676 33106 13688
rect 35618 13676 35624 13688
rect 35676 13676 35682 13728
rect 38194 13676 38200 13728
rect 38252 13676 38258 13728
rect 1104 13626 39192 13648
rect 1104 13574 5711 13626
rect 5763 13574 5775 13626
rect 5827 13574 5839 13626
rect 5891 13574 5903 13626
rect 5955 13574 5967 13626
rect 6019 13574 15233 13626
rect 15285 13574 15297 13626
rect 15349 13574 15361 13626
rect 15413 13574 15425 13626
rect 15477 13574 15489 13626
rect 15541 13574 24755 13626
rect 24807 13574 24819 13626
rect 24871 13574 24883 13626
rect 24935 13574 24947 13626
rect 24999 13574 25011 13626
rect 25063 13574 34277 13626
rect 34329 13574 34341 13626
rect 34393 13574 34405 13626
rect 34457 13574 34469 13626
rect 34521 13574 34533 13626
rect 34585 13574 39192 13626
rect 1104 13552 39192 13574
rect 3973 13515 4031 13521
rect 3973 13481 3985 13515
rect 4019 13512 4031 13515
rect 4062 13512 4068 13524
rect 4019 13484 4068 13512
rect 4019 13481 4031 13484
rect 3973 13475 4031 13481
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4172 13484 7236 13512
rect 2130 13404 2136 13456
rect 2188 13444 2194 13456
rect 2188 13416 2774 13444
rect 2188 13404 2194 13416
rect 2746 13376 2774 13416
rect 3694 13404 3700 13456
rect 3752 13444 3758 13456
rect 4172 13444 4200 13484
rect 3752 13416 4200 13444
rect 3752 13404 3758 13416
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 2746 13348 4537 13376
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 5442 13376 5448 13388
rect 4525 13339 4583 13345
rect 4632 13348 5448 13376
rect 1578 13268 1584 13320
rect 1636 13308 1642 13320
rect 2038 13308 2044 13320
rect 1636 13280 2044 13308
rect 1636 13268 1642 13280
rect 2038 13268 2044 13280
rect 2096 13308 2102 13320
rect 2593 13311 2651 13317
rect 2593 13308 2605 13311
rect 2096 13280 2605 13308
rect 2096 13268 2102 13280
rect 2593 13277 2605 13280
rect 2639 13308 2651 13311
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 2639 13280 3249 13308
rect 2639 13277 2651 13280
rect 2593 13271 2651 13277
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 3326 13268 3332 13320
rect 3384 13268 3390 13320
rect 4632 13308 4660 13348
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 5905 13379 5963 13385
rect 5905 13345 5917 13379
rect 5951 13376 5963 13379
rect 6546 13376 6552 13388
rect 5951 13348 6552 13376
rect 5951 13345 5963 13348
rect 5905 13339 5963 13345
rect 6546 13336 6552 13348
rect 6604 13376 6610 13388
rect 6914 13376 6920 13388
rect 6604 13348 6920 13376
rect 6604 13336 6610 13348
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 7208 13376 7236 13484
rect 7282 13472 7288 13524
rect 7340 13512 7346 13524
rect 8018 13512 8024 13524
rect 7340 13484 8024 13512
rect 7340 13472 7346 13484
rect 8018 13472 8024 13484
rect 8076 13512 8082 13524
rect 8297 13515 8355 13521
rect 8297 13512 8309 13515
rect 8076 13484 8309 13512
rect 8076 13472 8082 13484
rect 8297 13481 8309 13484
rect 8343 13481 8355 13515
rect 8297 13475 8355 13481
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 8527 13484 13019 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 7466 13404 7472 13456
rect 7524 13444 7530 13456
rect 12991 13444 13019 13484
rect 14274 13472 14280 13524
rect 14332 13512 14338 13524
rect 14550 13512 14556 13524
rect 14332 13484 14556 13512
rect 14332 13472 14338 13484
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 14734 13472 14740 13524
rect 14792 13472 14798 13524
rect 16025 13515 16083 13521
rect 16025 13481 16037 13515
rect 16071 13512 16083 13515
rect 16114 13512 16120 13524
rect 16071 13484 16120 13512
rect 16071 13481 16083 13484
rect 16025 13475 16083 13481
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 17126 13512 17132 13524
rect 16264 13484 17132 13512
rect 16264 13472 16270 13484
rect 17126 13472 17132 13484
rect 17184 13472 17190 13524
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 17770 13512 17776 13524
rect 17460 13484 17776 13512
rect 17460 13472 17466 13484
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 18414 13472 18420 13524
rect 18472 13472 18478 13524
rect 18782 13472 18788 13524
rect 18840 13472 18846 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 21140 13484 21772 13512
rect 21140 13472 21146 13484
rect 16301 13447 16359 13453
rect 16301 13444 16313 13447
rect 7524 13416 10916 13444
rect 12991 13416 16313 13444
rect 7524 13404 7530 13416
rect 7742 13376 7748 13388
rect 7208 13348 7748 13376
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 10781 13379 10839 13385
rect 10781 13376 10793 13379
rect 9824 13348 10793 13376
rect 9824 13336 9830 13348
rect 10781 13345 10793 13348
rect 10827 13345 10839 13379
rect 10888 13376 10916 13416
rect 16301 13413 16313 13416
rect 16347 13413 16359 13447
rect 16301 13407 16359 13413
rect 16574 13404 16580 13456
rect 16632 13444 16638 13456
rect 18279 13447 18337 13453
rect 18279 13444 18291 13447
rect 16632 13416 18291 13444
rect 16632 13404 16638 13416
rect 18279 13413 18291 13416
rect 18325 13413 18337 13447
rect 18279 13407 18337 13413
rect 19794 13404 19800 13456
rect 19852 13404 19858 13456
rect 21744 13444 21772 13484
rect 21818 13472 21824 13524
rect 21876 13512 21882 13524
rect 22830 13512 22836 13524
rect 21876 13484 22836 13512
rect 21876 13472 21882 13484
rect 22830 13472 22836 13484
rect 22888 13472 22894 13524
rect 23014 13472 23020 13524
rect 23072 13512 23078 13524
rect 23109 13515 23167 13521
rect 23109 13512 23121 13515
rect 23072 13484 23121 13512
rect 23072 13472 23078 13484
rect 23109 13481 23121 13484
rect 23155 13481 23167 13515
rect 23109 13475 23167 13481
rect 24949 13515 25007 13521
rect 24949 13481 24961 13515
rect 24995 13512 25007 13515
rect 32309 13515 32367 13521
rect 24995 13484 32260 13512
rect 24995 13481 25007 13484
rect 24949 13475 25007 13481
rect 23293 13447 23351 13453
rect 23293 13444 23305 13447
rect 21744 13416 23305 13444
rect 23293 13413 23305 13416
rect 23339 13413 23351 13447
rect 27341 13447 27399 13453
rect 27341 13444 27353 13447
rect 23293 13407 23351 13413
rect 24320 13416 27353 13444
rect 10888 13348 12296 13376
rect 10781 13339 10839 13345
rect 4080 13280 4660 13308
rect 1673 13243 1731 13249
rect 1673 13209 1685 13243
rect 1719 13240 1731 13243
rect 4080 13240 4108 13280
rect 5166 13268 5172 13320
rect 5224 13268 5230 13320
rect 9674 13268 9680 13320
rect 9732 13268 9738 13320
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 10321 13311 10379 13317
rect 10321 13308 10333 13311
rect 9916 13280 10333 13308
rect 9916 13268 9922 13280
rect 10321 13277 10333 13280
rect 10367 13277 10379 13311
rect 12268 13308 12296 13348
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 13262 13376 13268 13388
rect 12400 13348 13268 13376
rect 12400 13336 12406 13348
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13354 13336 13360 13388
rect 13412 13376 13418 13388
rect 13412 13348 13492 13376
rect 13412 13336 13418 13348
rect 12897 13311 12955 13317
rect 12268 13280 12434 13308
rect 10321 13271 10379 13277
rect 1719 13212 4108 13240
rect 4341 13243 4399 13249
rect 1719 13209 1731 13212
rect 1673 13203 1731 13209
rect 4341 13209 4353 13243
rect 4387 13240 4399 13243
rect 5350 13240 5356 13252
rect 4387 13212 5356 13240
rect 4387 13209 4399 13212
rect 4341 13203 4399 13209
rect 5350 13200 5356 13212
rect 5408 13200 5414 13252
rect 6178 13200 6184 13252
rect 6236 13200 6242 13252
rect 7834 13240 7840 13252
rect 7406 13212 7840 13240
rect 7834 13200 7840 13212
rect 7892 13200 7898 13252
rect 8113 13243 8171 13249
rect 8113 13209 8125 13243
rect 8159 13209 8171 13243
rect 8113 13203 8171 13209
rect 9769 13243 9827 13249
rect 9769 13209 9781 13243
rect 9815 13240 9827 13243
rect 9950 13240 9956 13252
rect 9815 13212 9956 13240
rect 9815 13209 9827 13212
rect 9769 13203 9827 13209
rect 934 13132 940 13184
rect 992 13172 998 13184
rect 1765 13175 1823 13181
rect 1765 13172 1777 13175
rect 992 13144 1777 13172
rect 992 13132 998 13144
rect 1765 13141 1777 13144
rect 1811 13141 1823 13175
rect 1765 13135 1823 13141
rect 2498 13132 2504 13184
rect 2556 13172 2562 13184
rect 2685 13175 2743 13181
rect 2685 13172 2697 13175
rect 2556 13144 2697 13172
rect 2556 13132 2562 13144
rect 2685 13141 2697 13144
rect 2731 13141 2743 13175
rect 2685 13135 2743 13141
rect 4430 13132 4436 13184
rect 4488 13132 4494 13184
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 5261 13175 5319 13181
rect 5261 13172 5273 13175
rect 4672 13144 5273 13172
rect 4672 13132 4678 13144
rect 5261 13141 5273 13144
rect 5307 13141 5319 13175
rect 5261 13135 5319 13141
rect 5994 13132 6000 13184
rect 6052 13172 6058 13184
rect 6362 13172 6368 13184
rect 6052 13144 6368 13172
rect 6052 13132 6058 13144
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 7653 13175 7711 13181
rect 7653 13141 7665 13175
rect 7699 13172 7711 13175
rect 8018 13172 8024 13184
rect 7699 13144 8024 13172
rect 7699 13141 7711 13144
rect 7653 13135 7711 13141
rect 8018 13132 8024 13144
rect 8076 13172 8082 13184
rect 8128 13172 8156 13203
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 10336 13212 11008 13240
rect 8076 13144 8156 13172
rect 8076 13132 8082 13144
rect 8294 13132 8300 13184
rect 8352 13181 8358 13184
rect 8352 13175 8371 13181
rect 8359 13141 8371 13175
rect 8352 13135 8371 13141
rect 8352 13132 8358 13135
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 10336 13172 10364 13212
rect 8812 13144 10364 13172
rect 10413 13175 10471 13181
rect 8812 13132 8818 13144
rect 10413 13141 10425 13175
rect 10459 13172 10471 13175
rect 10870 13172 10876 13184
rect 10459 13144 10876 13172
rect 10459 13141 10471 13144
rect 10413 13135 10471 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 10980 13172 11008 13212
rect 11054 13200 11060 13252
rect 11112 13200 11118 13252
rect 12066 13200 12072 13252
rect 12124 13200 12130 13252
rect 12406 13240 12434 13280
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 13170 13308 13176 13320
rect 12943 13280 13176 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 13464 13317 13492 13348
rect 13556 13348 15056 13376
rect 13556 13317 13584 13348
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 14918 13308 14924 13320
rect 13688 13280 14924 13308
rect 13688 13268 13694 13280
rect 14918 13268 14924 13280
rect 14976 13268 14982 13320
rect 15028 13308 15056 13348
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 15252 13348 15301 13376
rect 15252 13336 15258 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 15289 13339 15347 13345
rect 16022 13336 16028 13388
rect 16080 13376 16086 13388
rect 16666 13376 16672 13388
rect 16080 13348 16672 13376
rect 16080 13336 16086 13348
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 18509 13379 18567 13385
rect 18509 13376 18521 13379
rect 16908 13348 18521 13376
rect 16908 13336 16914 13348
rect 18509 13345 18521 13348
rect 18555 13345 18567 13379
rect 18509 13339 18567 13345
rect 15746 13308 15752 13320
rect 15028 13280 15752 13308
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 16114 13268 16120 13320
rect 16172 13308 16178 13320
rect 16393 13311 16451 13317
rect 16393 13308 16405 13311
rect 16172 13280 16405 13308
rect 16172 13268 16178 13280
rect 16393 13277 16405 13280
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13277 16543 13311
rect 16485 13271 16543 13277
rect 12406 13212 13124 13240
rect 12342 13172 12348 13184
rect 10980 13144 12348 13172
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12529 13175 12587 13181
rect 12529 13172 12541 13175
rect 12492 13144 12541 13172
rect 12492 13132 12498 13144
rect 12529 13141 12541 13144
rect 12575 13141 12587 13175
rect 13096 13172 13124 13212
rect 13262 13200 13268 13252
rect 13320 13240 13326 13252
rect 13357 13243 13415 13249
rect 13357 13240 13369 13243
rect 13320 13212 13369 13240
rect 13320 13200 13326 13212
rect 13357 13209 13369 13212
rect 13403 13240 13415 13243
rect 13403 13212 14228 13240
rect 13403 13209 13415 13212
rect 13357 13203 13415 13209
rect 13725 13175 13783 13181
rect 13725 13172 13737 13175
rect 13096 13144 13737 13172
rect 12529 13135 12587 13141
rect 13725 13141 13737 13144
rect 13771 13141 13783 13175
rect 14200 13172 14228 13212
rect 14274 13200 14280 13252
rect 14332 13240 14338 13252
rect 15197 13243 15255 13249
rect 15197 13240 15209 13243
rect 14332 13212 15209 13240
rect 14332 13200 14338 13212
rect 15197 13209 15209 13212
rect 15243 13240 15255 13243
rect 15654 13240 15660 13252
rect 15243 13212 15660 13240
rect 15243 13209 15255 13212
rect 15197 13203 15255 13209
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 16500 13240 16528 13271
rect 16758 13268 16764 13320
rect 16816 13268 16822 13320
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13308 17279 13311
rect 18690 13308 18696 13320
rect 17267 13280 18696 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 19426 13268 19432 13320
rect 19484 13268 19490 13320
rect 19518 13268 19524 13320
rect 19576 13308 19582 13320
rect 19812 13317 19840 13404
rect 20441 13379 20499 13385
rect 20441 13345 20453 13379
rect 20487 13376 20499 13379
rect 20714 13376 20720 13388
rect 20487 13348 20720 13376
rect 20487 13345 20499 13348
rect 20441 13339 20499 13345
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 21266 13336 21272 13388
rect 21324 13376 21330 13388
rect 24320 13376 24348 13416
rect 27341 13413 27353 13416
rect 27387 13413 27399 13447
rect 27341 13407 27399 13413
rect 27430 13404 27436 13456
rect 27488 13444 27494 13456
rect 27488 13416 28580 13444
rect 27488 13404 27494 13416
rect 21324 13348 24348 13376
rect 25593 13379 25651 13385
rect 21324 13336 21330 13348
rect 25593 13345 25605 13379
rect 25639 13376 25651 13379
rect 26142 13376 26148 13388
rect 25639 13348 26148 13376
rect 25639 13345 25651 13348
rect 25593 13339 25651 13345
rect 26142 13336 26148 13348
rect 26200 13336 26206 13388
rect 26602 13336 26608 13388
rect 26660 13336 26666 13388
rect 26789 13379 26847 13385
rect 26789 13345 26801 13379
rect 26835 13376 26847 13379
rect 27706 13376 27712 13388
rect 26835 13348 27712 13376
rect 26835 13345 26847 13348
rect 26789 13339 26847 13345
rect 27706 13336 27712 13348
rect 27764 13336 27770 13388
rect 27982 13336 27988 13388
rect 28040 13336 28046 13388
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19576 13280 19625 13308
rect 19576 13268 19582 13280
rect 19613 13277 19625 13280
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 22186 13268 22192 13320
rect 22244 13308 22250 13320
rect 22370 13308 22376 13320
rect 22244 13280 22376 13308
rect 22244 13268 22250 13280
rect 22370 13268 22376 13280
rect 22428 13268 22434 13320
rect 22465 13311 22523 13317
rect 22465 13277 22477 13311
rect 22511 13308 22523 13311
rect 22738 13308 22744 13320
rect 22511 13280 22744 13308
rect 22511 13277 22523 13280
rect 22465 13271 22523 13277
rect 22738 13268 22744 13280
rect 22796 13268 22802 13320
rect 22830 13268 22836 13320
rect 22888 13308 22894 13320
rect 22888 13280 23428 13308
rect 22888 13268 22894 13280
rect 16942 13240 16948 13252
rect 16500 13212 16948 13240
rect 16942 13200 16948 13212
rect 17000 13200 17006 13252
rect 17497 13243 17555 13249
rect 17497 13209 17509 13243
rect 17543 13240 17555 13243
rect 17678 13240 17684 13252
rect 17543 13212 17684 13240
rect 17543 13209 17555 13212
rect 17497 13203 17555 13209
rect 17678 13200 17684 13212
rect 17736 13200 17742 13252
rect 18138 13200 18144 13252
rect 18196 13200 18202 13252
rect 18230 13200 18236 13252
rect 18288 13240 18294 13252
rect 18414 13240 18420 13252
rect 18288 13212 18420 13240
rect 18288 13200 18294 13212
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 19705 13243 19763 13249
rect 19705 13209 19717 13243
rect 19751 13240 19763 13243
rect 20438 13240 20444 13252
rect 19751 13212 20444 13240
rect 19751 13209 19763 13212
rect 19705 13203 19763 13209
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 20717 13243 20775 13249
rect 20717 13209 20729 13243
rect 20763 13209 20775 13243
rect 22002 13240 22008 13252
rect 21942 13212 22008 13240
rect 20717 13203 20775 13209
rect 14734 13172 14740 13184
rect 14200 13144 14740 13172
rect 13725 13135 13783 13141
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 14918 13132 14924 13184
rect 14976 13172 14982 13184
rect 15105 13175 15163 13181
rect 15105 13172 15117 13175
rect 14976 13144 15117 13172
rect 14976 13132 14982 13144
rect 15105 13141 15117 13144
rect 15151 13141 15163 13175
rect 15105 13135 15163 13141
rect 15286 13132 15292 13184
rect 15344 13172 15350 13184
rect 16669 13175 16727 13181
rect 16669 13172 16681 13175
rect 15344 13144 16681 13172
rect 15344 13132 15350 13144
rect 16669 13141 16681 13144
rect 16715 13141 16727 13175
rect 16669 13135 16727 13141
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 19886 13172 19892 13184
rect 16816 13144 19892 13172
rect 16816 13132 16822 13144
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 19981 13175 20039 13181
rect 19981 13141 19993 13175
rect 20027 13172 20039 13175
rect 20346 13172 20352 13184
rect 20027 13144 20352 13172
rect 20027 13141 20039 13144
rect 19981 13135 20039 13141
rect 20346 13132 20352 13144
rect 20404 13132 20410 13184
rect 20732 13172 20760 13203
rect 22002 13200 22008 13212
rect 22060 13200 22066 13252
rect 22554 13240 22560 13252
rect 22112 13212 22560 13240
rect 22112 13172 22140 13212
rect 22554 13200 22560 13212
rect 22612 13200 22618 13252
rect 22925 13243 22983 13249
rect 22925 13209 22937 13243
rect 22971 13240 22983 13243
rect 23290 13240 23296 13252
rect 22971 13212 23296 13240
rect 22971 13209 22983 13212
rect 22925 13203 22983 13209
rect 23290 13200 23296 13212
rect 23348 13200 23354 13252
rect 23400 13240 23428 13280
rect 23842 13268 23848 13320
rect 23900 13268 23906 13320
rect 24578 13268 24584 13320
rect 24636 13308 24642 13320
rect 28552 13317 28580 13416
rect 28902 13404 28908 13456
rect 28960 13444 28966 13456
rect 30282 13444 30288 13456
rect 28960 13416 30288 13444
rect 28960 13404 28966 13416
rect 30282 13404 30288 13416
rect 30340 13404 30346 13456
rect 32232 13444 32260 13484
rect 32309 13481 32321 13515
rect 32355 13512 32367 13515
rect 32766 13512 32772 13524
rect 32355 13484 32772 13512
rect 32355 13481 32367 13484
rect 32309 13475 32367 13481
rect 32766 13472 32772 13484
rect 32824 13512 32830 13524
rect 33042 13512 33048 13524
rect 32824 13484 33048 13512
rect 32824 13472 32830 13484
rect 33042 13472 33048 13484
rect 33100 13472 33106 13524
rect 33686 13472 33692 13524
rect 33744 13512 33750 13524
rect 36633 13515 36691 13521
rect 36633 13512 36645 13515
rect 33744 13484 36645 13512
rect 33744 13472 33750 13484
rect 36633 13481 36645 13484
rect 36679 13481 36691 13515
rect 36633 13475 36691 13481
rect 33962 13444 33968 13456
rect 32232 13416 33968 13444
rect 33962 13404 33968 13416
rect 34020 13404 34026 13456
rect 34054 13404 34060 13456
rect 34112 13404 34118 13456
rect 29914 13336 29920 13388
rect 29972 13376 29978 13388
rect 30561 13379 30619 13385
rect 30561 13376 30573 13379
rect 29972 13348 30573 13376
rect 29972 13336 29978 13348
rect 30561 13345 30573 13348
rect 30607 13376 30619 13379
rect 30926 13376 30932 13388
rect 30607 13348 30932 13376
rect 30607 13345 30619 13348
rect 30561 13339 30619 13345
rect 30926 13336 30932 13348
rect 30984 13336 30990 13388
rect 32398 13336 32404 13388
rect 32456 13376 32462 13388
rect 33321 13379 33379 13385
rect 33321 13376 33333 13379
rect 32456 13348 33333 13376
rect 32456 13336 32462 13348
rect 33321 13345 33333 13348
rect 33367 13376 33379 13379
rect 34790 13376 34796 13388
rect 33367 13348 34796 13376
rect 33367 13345 33379 13348
rect 33321 13339 33379 13345
rect 34790 13336 34796 13348
rect 34848 13336 34854 13388
rect 34882 13336 34888 13388
rect 34940 13336 34946 13388
rect 25409 13311 25467 13317
rect 25409 13308 25421 13311
rect 24636 13280 25421 13308
rect 24636 13268 24642 13280
rect 25409 13277 25421 13280
rect 25455 13277 25467 13311
rect 27801 13311 27859 13317
rect 27801 13308 27813 13311
rect 25409 13271 25467 13277
rect 25700 13280 27813 13308
rect 25317 13243 25375 13249
rect 23400 13212 24072 13240
rect 20732 13144 22140 13172
rect 22186 13132 22192 13184
rect 22244 13172 22250 13184
rect 23125 13175 23183 13181
rect 23125 13172 23137 13175
rect 22244 13144 23137 13172
rect 22244 13132 22250 13144
rect 23125 13141 23137 13144
rect 23171 13172 23183 13175
rect 23658 13172 23664 13184
rect 23171 13144 23664 13172
rect 23171 13141 23183 13144
rect 23125 13135 23183 13141
rect 23658 13132 23664 13144
rect 23716 13132 23722 13184
rect 23934 13132 23940 13184
rect 23992 13132 23998 13184
rect 24044 13172 24072 13212
rect 25317 13209 25329 13243
rect 25363 13240 25375 13243
rect 25590 13240 25596 13252
rect 25363 13212 25596 13240
rect 25363 13209 25375 13212
rect 25317 13203 25375 13209
rect 25590 13200 25596 13212
rect 25648 13200 25654 13252
rect 25700 13172 25728 13280
rect 27801 13277 27813 13280
rect 27847 13277 27859 13311
rect 27801 13271 27859 13277
rect 28537 13311 28595 13317
rect 28537 13277 28549 13311
rect 28583 13308 28595 13311
rect 29733 13311 29791 13317
rect 29733 13308 29745 13311
rect 28583 13280 29745 13308
rect 28583 13277 28595 13280
rect 28537 13271 28595 13277
rect 29733 13277 29745 13280
rect 29779 13308 29791 13311
rect 30190 13308 30196 13320
rect 29779 13280 30196 13308
rect 29779 13277 29791 13280
rect 29733 13271 29791 13277
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 33137 13311 33195 13317
rect 33137 13277 33149 13311
rect 33183 13308 33195 13311
rect 33686 13308 33692 13320
rect 33183 13280 33692 13308
rect 33183 13277 33195 13280
rect 33137 13271 33195 13277
rect 33686 13268 33692 13280
rect 33744 13268 33750 13320
rect 33870 13268 33876 13320
rect 33928 13308 33934 13320
rect 33965 13311 34023 13317
rect 33965 13308 33977 13311
rect 33928 13280 33977 13308
rect 33928 13268 33934 13280
rect 33965 13277 33977 13280
rect 34011 13277 34023 13311
rect 33965 13271 34023 13277
rect 37553 13311 37611 13317
rect 37553 13277 37565 13311
rect 37599 13308 37611 13311
rect 38378 13308 38384 13320
rect 37599 13280 38384 13308
rect 37599 13277 37611 13280
rect 37553 13271 37611 13277
rect 38378 13268 38384 13280
rect 38436 13268 38442 13320
rect 26786 13200 26792 13252
rect 26844 13240 26850 13252
rect 27709 13243 27767 13249
rect 27709 13240 27721 13243
rect 26844 13212 27721 13240
rect 26844 13200 26850 13212
rect 27709 13209 27721 13212
rect 27755 13209 27767 13243
rect 27709 13203 27767 13209
rect 28166 13200 28172 13252
rect 28224 13240 28230 13252
rect 29825 13243 29883 13249
rect 29825 13240 29837 13243
rect 28224 13212 29837 13240
rect 28224 13200 28230 13212
rect 29825 13209 29837 13212
rect 29871 13209 29883 13243
rect 29825 13203 29883 13209
rect 30834 13200 30840 13252
rect 30892 13200 30898 13252
rect 31846 13200 31852 13252
rect 31904 13200 31910 13252
rect 35161 13243 35219 13249
rect 35161 13240 35173 13243
rect 32784 13212 35173 13240
rect 24044 13144 25728 13172
rect 25866 13132 25872 13184
rect 25924 13172 25930 13184
rect 26145 13175 26203 13181
rect 26145 13172 26157 13175
rect 25924 13144 26157 13172
rect 25924 13132 25930 13144
rect 26145 13141 26157 13144
rect 26191 13141 26203 13175
rect 26145 13135 26203 13141
rect 26510 13132 26516 13184
rect 26568 13132 26574 13184
rect 28442 13132 28448 13184
rect 28500 13172 28506 13184
rect 28629 13175 28687 13181
rect 28629 13172 28641 13175
rect 28500 13144 28641 13172
rect 28500 13132 28506 13144
rect 28629 13141 28641 13144
rect 28675 13141 28687 13175
rect 28629 13135 28687 13141
rect 28810 13132 28816 13184
rect 28868 13172 28874 13184
rect 30466 13172 30472 13184
rect 28868 13144 30472 13172
rect 28868 13132 28874 13144
rect 30466 13132 30472 13144
rect 30524 13132 30530 13184
rect 32784 13181 32812 13212
rect 35161 13209 35173 13212
rect 35207 13209 35219 13243
rect 38194 13240 38200 13252
rect 36386 13212 38200 13240
rect 35161 13203 35219 13209
rect 38194 13200 38200 13212
rect 38252 13200 38258 13252
rect 38289 13243 38347 13249
rect 38289 13209 38301 13243
rect 38335 13240 38347 13243
rect 39390 13240 39396 13252
rect 38335 13212 39396 13240
rect 38335 13209 38347 13212
rect 38289 13203 38347 13209
rect 39390 13200 39396 13212
rect 39448 13200 39454 13252
rect 32769 13175 32827 13181
rect 32769 13141 32781 13175
rect 32815 13141 32827 13175
rect 32769 13135 32827 13141
rect 32858 13132 32864 13184
rect 32916 13172 32922 13184
rect 33229 13175 33287 13181
rect 33229 13172 33241 13175
rect 32916 13144 33241 13172
rect 32916 13132 32922 13144
rect 33229 13141 33241 13144
rect 33275 13172 33287 13175
rect 35894 13172 35900 13184
rect 33275 13144 35900 13172
rect 33275 13141 33287 13144
rect 33229 13135 33287 13141
rect 35894 13132 35900 13144
rect 35952 13132 35958 13184
rect 37366 13132 37372 13184
rect 37424 13172 37430 13184
rect 37645 13175 37703 13181
rect 37645 13172 37657 13175
rect 37424 13144 37657 13172
rect 37424 13132 37430 13144
rect 37645 13141 37657 13144
rect 37691 13141 37703 13175
rect 37645 13135 37703 13141
rect 37734 13132 37740 13184
rect 37792 13172 37798 13184
rect 38381 13175 38439 13181
rect 38381 13172 38393 13175
rect 37792 13144 38393 13172
rect 37792 13132 37798 13144
rect 38381 13141 38393 13144
rect 38427 13141 38439 13175
rect 38381 13135 38439 13141
rect 1104 13082 39352 13104
rect 1104 13030 10472 13082
rect 10524 13030 10536 13082
rect 10588 13030 10600 13082
rect 10652 13030 10664 13082
rect 10716 13030 10728 13082
rect 10780 13030 19994 13082
rect 20046 13030 20058 13082
rect 20110 13030 20122 13082
rect 20174 13030 20186 13082
rect 20238 13030 20250 13082
rect 20302 13030 29516 13082
rect 29568 13030 29580 13082
rect 29632 13030 29644 13082
rect 29696 13030 29708 13082
rect 29760 13030 29772 13082
rect 29824 13030 39038 13082
rect 39090 13030 39102 13082
rect 39154 13030 39166 13082
rect 39218 13030 39230 13082
rect 39282 13030 39294 13082
rect 39346 13030 39352 13082
rect 1104 13008 39352 13030
rect 6086 12968 6092 12980
rect 2516 12940 6092 12968
rect 2516 12909 2544 12940
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 7561 12971 7619 12977
rect 7561 12968 7573 12971
rect 6236 12940 7573 12968
rect 6236 12928 6242 12940
rect 7561 12937 7573 12940
rect 7607 12937 7619 12971
rect 7561 12931 7619 12937
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7800 12940 7941 12968
rect 7800 12928 7806 12940
rect 7929 12937 7941 12940
rect 7975 12937 7987 12971
rect 7929 12931 7987 12937
rect 8018 12928 8024 12980
rect 8076 12928 8082 12980
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 8352 12940 11008 12968
rect 8352 12928 8358 12940
rect 2501 12903 2559 12909
rect 2501 12869 2513 12903
rect 2547 12869 2559 12903
rect 2501 12863 2559 12869
rect 3510 12860 3516 12912
rect 3568 12860 3574 12912
rect 3786 12860 3792 12912
rect 3844 12900 3850 12912
rect 4249 12903 4307 12909
rect 4249 12900 4261 12903
rect 3844 12872 4261 12900
rect 3844 12860 3850 12872
rect 4249 12869 4261 12872
rect 4295 12869 4307 12903
rect 4249 12863 4307 12869
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 4488 12872 7696 12900
rect 4488 12860 4494 12872
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 2038 12832 2044 12844
rect 1627 12804 2044 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 5166 12832 5172 12844
rect 4908 12804 5172 12832
rect 2222 12724 2228 12776
rect 2280 12724 2286 12776
rect 4522 12764 4528 12776
rect 2332 12736 4528 12764
rect 1946 12656 1952 12708
rect 2004 12696 2010 12708
rect 2332 12696 2360 12736
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 2004 12668 2360 12696
rect 2004 12656 2010 12668
rect 3602 12656 3608 12708
rect 3660 12696 3666 12708
rect 4908 12696 4936 12804
rect 5166 12792 5172 12804
rect 5224 12832 5230 12844
rect 5626 12832 5632 12844
rect 5224 12804 5632 12832
rect 5224 12792 5230 12804
rect 5626 12792 5632 12804
rect 5684 12832 5690 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5684 12804 5825 12832
rect 5684 12792 5690 12804
rect 5813 12801 5825 12804
rect 5859 12832 5871 12835
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 5859 12804 6929 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6917 12801 6929 12804
rect 6963 12832 6975 12835
rect 7558 12832 7564 12844
rect 6963 12804 7564 12832
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 7668 12832 7696 12872
rect 7834 12860 7840 12912
rect 7892 12900 7898 12912
rect 9769 12903 9827 12909
rect 9769 12900 9781 12903
rect 7892 12872 9781 12900
rect 7892 12860 7898 12872
rect 9769 12869 9781 12872
rect 9815 12869 9827 12903
rect 10980 12900 11008 12940
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11701 12971 11759 12977
rect 11701 12968 11713 12971
rect 11112 12940 11713 12968
rect 11112 12928 11118 12940
rect 11701 12937 11713 12940
rect 11747 12937 11759 12971
rect 11701 12931 11759 12937
rect 13096 12940 13492 12968
rect 13096 12900 13124 12940
rect 10980 12872 13124 12900
rect 9769 12863 9827 12869
rect 13170 12860 13176 12912
rect 13228 12860 13234 12912
rect 13262 12860 13268 12912
rect 13320 12900 13326 12912
rect 13373 12903 13431 12909
rect 13373 12900 13385 12903
rect 13320 12872 13385 12900
rect 13320 12860 13326 12872
rect 13373 12869 13385 12872
rect 13419 12869 13431 12903
rect 13464 12900 13492 12940
rect 13538 12928 13544 12980
rect 13596 12928 13602 12980
rect 13648 12940 14596 12968
rect 13648 12900 13676 12940
rect 13464 12872 13676 12900
rect 14568 12900 14596 12940
rect 14642 12928 14648 12980
rect 14700 12968 14706 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 14700 12940 14749 12968
rect 14700 12928 14706 12940
rect 14737 12937 14749 12940
rect 14783 12937 14795 12971
rect 14737 12931 14795 12937
rect 14918 12928 14924 12980
rect 14976 12968 14982 12980
rect 15194 12968 15200 12980
rect 14976 12940 15200 12968
rect 14976 12928 14982 12940
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 16133 12971 16191 12977
rect 16133 12968 16145 12971
rect 15304 12940 16145 12968
rect 15304 12900 15332 12940
rect 16133 12937 16145 12940
rect 16179 12968 16191 12971
rect 16390 12968 16396 12980
rect 16179 12940 16396 12968
rect 16179 12937 16191 12940
rect 16133 12931 16191 12937
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 16482 12928 16488 12980
rect 16540 12968 16546 12980
rect 16540 12940 16712 12968
rect 16540 12928 16546 12940
rect 15959 12903 16017 12909
rect 15959 12900 15971 12903
rect 14568 12872 15332 12900
rect 13373 12863 13431 12869
rect 15948 12869 15971 12900
rect 16005 12869 16017 12903
rect 16684 12900 16712 12940
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 18601 12971 18659 12977
rect 18601 12968 18613 12971
rect 16816 12940 18613 12968
rect 16816 12928 16822 12940
rect 18601 12937 18613 12940
rect 18647 12937 18659 12971
rect 18601 12931 18659 12937
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 18874 12968 18880 12980
rect 18748 12940 18880 12968
rect 18748 12928 18754 12940
rect 18874 12928 18880 12940
rect 18932 12928 18938 12980
rect 20714 12968 20720 12980
rect 19076 12940 20720 12968
rect 17129 12903 17187 12909
rect 17129 12900 17141 12903
rect 15948 12863 16017 12869
rect 16224 12872 16436 12900
rect 16684 12872 17141 12900
rect 7668 12804 8340 12832
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 5951 12736 7420 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 7190 12696 7196 12708
rect 3660 12668 4936 12696
rect 5000 12668 7196 12696
rect 3660 12656 3666 12668
rect 1673 12631 1731 12637
rect 1673 12597 1685 12631
rect 1719 12628 1731 12631
rect 5000 12628 5028 12668
rect 7190 12656 7196 12668
rect 7248 12656 7254 12708
rect 7392 12696 7420 12736
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 8202 12764 8208 12776
rect 7524 12736 8208 12764
rect 7524 12724 7530 12736
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8312 12764 8340 12804
rect 8754 12792 8760 12844
rect 8812 12792 8818 12844
rect 8864 12804 9076 12832
rect 8864 12764 8892 12804
rect 8312 12736 8892 12764
rect 8938 12724 8944 12776
rect 8996 12724 9002 12776
rect 9048 12764 9076 12804
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 9950 12832 9956 12844
rect 9732 12804 9956 12832
rect 9732 12792 9738 12804
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 10192 12804 10333 12832
rect 10192 12792 10198 12804
rect 10321 12801 10333 12804
rect 10367 12832 10379 12835
rect 10502 12832 10508 12844
rect 10367 12804 10508 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 10502 12792 10508 12804
rect 10560 12832 10566 12844
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10560 12804 10977 12832
rect 10560 12792 10566 12804
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 12066 12792 12072 12844
rect 12124 12792 12130 12844
rect 12158 12792 12164 12844
rect 12216 12832 12222 12844
rect 12894 12832 12900 12844
rect 12216 12830 12296 12832
rect 12452 12830 12900 12832
rect 12216 12804 12900 12830
rect 12216 12792 12222 12804
rect 12268 12802 12480 12804
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14001 12835 14059 12841
rect 14001 12832 14013 12835
rect 13872 12804 14013 12832
rect 13872 12792 13878 12804
rect 14001 12801 14013 12804
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12832 14151 12835
rect 15102 12832 15108 12844
rect 14139 12804 15108 12832
rect 14139 12801 14151 12804
rect 14093 12795 14151 12801
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15654 12832 15660 12844
rect 15335 12804 15660 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 15838 12792 15844 12844
rect 15896 12832 15902 12844
rect 15948 12832 15976 12863
rect 15896 12804 15976 12832
rect 15896 12792 15902 12804
rect 10870 12764 10876 12776
rect 9048 12736 10876 12764
rect 10870 12724 10876 12736
rect 10928 12724 10934 12776
rect 12345 12767 12403 12773
rect 12345 12764 12357 12767
rect 12268 12736 12357 12764
rect 12268 12708 12296 12736
rect 12345 12733 12357 12736
rect 12391 12733 12403 12767
rect 12345 12727 12403 12733
rect 13722 12724 13728 12776
rect 13780 12764 13786 12776
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 13780 12736 15209 12764
rect 13780 12724 13786 12736
rect 15197 12733 15209 12736
rect 15243 12733 15255 12767
rect 15197 12727 15255 12733
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12764 15531 12767
rect 15746 12764 15752 12776
rect 15519 12736 15752 12764
rect 15519 12733 15531 12736
rect 15473 12727 15531 12733
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 15930 12724 15936 12776
rect 15988 12764 15994 12776
rect 16224 12764 16252 12872
rect 16408 12832 16436 12872
rect 17129 12869 17141 12872
rect 17175 12869 17187 12903
rect 18966 12900 18972 12912
rect 18354 12872 18972 12900
rect 17129 12863 17187 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 19076 12841 19104 12940
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 25225 12971 25283 12977
rect 25225 12968 25237 12971
rect 22066 12940 25237 12968
rect 22066 12900 22094 12940
rect 25225 12937 25237 12940
rect 25271 12937 25283 12971
rect 25225 12931 25283 12937
rect 25498 12928 25504 12980
rect 25556 12968 25562 12980
rect 25869 12971 25927 12977
rect 25869 12968 25881 12971
rect 25556 12940 25881 12968
rect 25556 12928 25562 12940
rect 25869 12937 25881 12940
rect 25915 12937 25927 12971
rect 25869 12931 25927 12937
rect 26234 12928 26240 12980
rect 26292 12968 26298 12980
rect 26329 12971 26387 12977
rect 26329 12968 26341 12971
rect 26292 12940 26341 12968
rect 26292 12928 26298 12940
rect 26329 12937 26341 12940
rect 26375 12937 26387 12971
rect 26329 12931 26387 12937
rect 26510 12928 26516 12980
rect 26568 12968 26574 12980
rect 26568 12940 29040 12968
rect 26568 12928 26574 12940
rect 22830 12900 22836 12912
rect 20562 12872 22094 12900
rect 22204 12872 22836 12900
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16408 12804 16865 12832
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12801 19119 12835
rect 21266 12832 21272 12844
rect 19061 12795 19119 12801
rect 21008 12804 21272 12832
rect 15988 12736 16252 12764
rect 19337 12767 19395 12773
rect 15988 12724 15994 12736
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 21008 12764 21036 12804
rect 21266 12792 21272 12804
rect 21324 12792 21330 12844
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21968 12804 22017 12832
rect 21968 12792 21974 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22204 12832 22232 12872
rect 22830 12860 22836 12872
rect 22888 12860 22894 12912
rect 23106 12860 23112 12912
rect 23164 12900 23170 12912
rect 23164 12872 23690 12900
rect 23164 12860 23170 12872
rect 26142 12860 26148 12912
rect 26200 12900 26206 12912
rect 27982 12900 27988 12912
rect 26200 12872 27988 12900
rect 26200 12860 26206 12872
rect 27982 12860 27988 12872
rect 28040 12900 28046 12912
rect 28350 12900 28356 12912
rect 28040 12872 28356 12900
rect 28040 12860 28046 12872
rect 28350 12860 28356 12872
rect 28408 12860 28414 12912
rect 29012 12909 29040 12940
rect 31478 12928 31484 12980
rect 31536 12928 31542 12980
rect 31754 12928 31760 12980
rect 31812 12968 31818 12980
rect 32858 12968 32864 12980
rect 31812 12940 32864 12968
rect 31812 12928 31818 12940
rect 32858 12928 32864 12940
rect 32916 12928 32922 12980
rect 33134 12928 33140 12980
rect 33192 12968 33198 12980
rect 33410 12968 33416 12980
rect 33192 12940 33416 12968
rect 33192 12928 33198 12940
rect 33410 12928 33416 12940
rect 33468 12928 33474 12980
rect 35250 12968 35256 12980
rect 33520 12940 35256 12968
rect 28905 12903 28963 12909
rect 28905 12900 28917 12903
rect 28460 12872 28917 12900
rect 22005 12795 22063 12801
rect 22112 12804 22232 12832
rect 19383 12736 21036 12764
rect 21085 12767 21143 12773
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 21085 12733 21097 12767
rect 21131 12764 21143 12767
rect 22112 12764 22140 12804
rect 22370 12792 22376 12844
rect 22428 12832 22434 12844
rect 22922 12832 22928 12844
rect 22428 12804 22928 12832
rect 22428 12792 22434 12804
rect 22922 12792 22928 12804
rect 22980 12792 22986 12844
rect 24486 12792 24492 12844
rect 24544 12832 24550 12844
rect 25133 12835 25191 12841
rect 25133 12832 25145 12835
rect 24544 12804 25145 12832
rect 24544 12792 24550 12804
rect 25133 12801 25145 12804
rect 25179 12832 25191 12835
rect 25866 12832 25872 12844
rect 25179 12804 25872 12832
rect 25179 12801 25191 12804
rect 25133 12795 25191 12801
rect 25866 12792 25872 12804
rect 25924 12792 25930 12844
rect 26234 12792 26240 12844
rect 26292 12792 26298 12844
rect 27525 12835 27583 12841
rect 27525 12801 27537 12835
rect 27571 12832 27583 12835
rect 28074 12832 28080 12844
rect 27571 12804 28080 12832
rect 27571 12801 27583 12804
rect 27525 12795 27583 12801
rect 28074 12792 28080 12804
rect 28132 12792 28138 12844
rect 28258 12792 28264 12844
rect 28316 12832 28322 12844
rect 28460 12832 28488 12872
rect 28905 12869 28917 12872
rect 28951 12869 28963 12903
rect 28905 12863 28963 12869
rect 28997 12903 29055 12909
rect 28997 12869 29009 12903
rect 29043 12869 29055 12903
rect 29914 12900 29920 12912
rect 28997 12863 29055 12869
rect 29748 12872 29920 12900
rect 28316 12804 28488 12832
rect 28316 12792 28322 12804
rect 28718 12792 28724 12844
rect 28776 12792 28782 12844
rect 29086 12792 29092 12844
rect 29144 12792 29150 12844
rect 29362 12792 29368 12844
rect 29420 12832 29426 12844
rect 29748 12841 29776 12872
rect 29914 12860 29920 12872
rect 29972 12860 29978 12912
rect 30006 12860 30012 12912
rect 30064 12860 30070 12912
rect 32674 12860 32680 12912
rect 32732 12900 32738 12912
rect 32953 12903 33011 12909
rect 32953 12900 32965 12903
rect 32732 12872 32965 12900
rect 32732 12860 32738 12872
rect 32953 12869 32965 12872
rect 32999 12869 33011 12903
rect 33520 12900 33548 12940
rect 35250 12928 35256 12940
rect 35308 12968 35314 12980
rect 35434 12968 35440 12980
rect 35308 12940 35440 12968
rect 35308 12928 35314 12940
rect 35434 12928 35440 12940
rect 35492 12928 35498 12980
rect 32953 12863 33011 12869
rect 33152 12872 33548 12900
rect 34885 12903 34943 12909
rect 29733 12835 29791 12841
rect 29733 12832 29745 12835
rect 29420 12804 29745 12832
rect 29420 12792 29426 12804
rect 29733 12801 29745 12804
rect 29779 12801 29791 12835
rect 32769 12835 32827 12841
rect 31142 12804 31892 12832
rect 29733 12795 29791 12801
rect 21131 12736 22140 12764
rect 21131 12733 21143 12736
rect 21085 12727 21143 12733
rect 22186 12724 22192 12776
rect 22244 12724 22250 12776
rect 23201 12767 23259 12773
rect 23201 12764 23213 12767
rect 22388 12736 23213 12764
rect 22388 12708 22416 12736
rect 23201 12733 23213 12736
rect 23247 12733 23259 12767
rect 23201 12727 23259 12733
rect 26513 12767 26571 12773
rect 26513 12733 26525 12767
rect 26559 12764 26571 12767
rect 26602 12764 26608 12776
rect 26559 12736 26608 12764
rect 26559 12733 26571 12736
rect 26513 12727 26571 12733
rect 26602 12724 26608 12736
rect 26660 12764 26666 12776
rect 28810 12764 28816 12776
rect 26660 12736 28816 12764
rect 26660 12724 26666 12736
rect 28810 12724 28816 12736
rect 28868 12724 28874 12776
rect 31754 12764 31760 12776
rect 29840 12736 31760 12764
rect 7392 12668 9628 12696
rect 1719 12600 5028 12628
rect 1719 12597 1731 12600
rect 1673 12591 1731 12597
rect 5258 12588 5264 12640
rect 5316 12588 5322 12640
rect 7009 12631 7067 12637
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 9214 12628 9220 12640
rect 7055 12600 9220 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 9600 12628 9628 12668
rect 9674 12656 9680 12708
rect 9732 12696 9738 12708
rect 10413 12699 10471 12705
rect 9732 12668 10272 12696
rect 9732 12656 9738 12668
rect 10134 12628 10140 12640
rect 9600 12600 10140 12628
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 10244 12628 10272 12668
rect 10413 12665 10425 12699
rect 10459 12696 10471 12699
rect 11514 12696 11520 12708
rect 10459 12668 11520 12696
rect 10459 12665 10471 12668
rect 10413 12659 10471 12665
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 12250 12656 12256 12708
rect 12308 12696 12314 12708
rect 14642 12696 14648 12708
rect 12308 12668 14648 12696
rect 12308 12656 12314 12668
rect 14642 12656 14648 12668
rect 14700 12656 14706 12708
rect 15013 12699 15071 12705
rect 15013 12665 15025 12699
rect 15059 12696 15071 12699
rect 16301 12699 16359 12705
rect 16301 12696 16313 12699
rect 15059 12668 15608 12696
rect 15059 12665 15071 12668
rect 15013 12659 15071 12665
rect 10778 12628 10784 12640
rect 10244 12600 10784 12628
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11057 12631 11115 12637
rect 11057 12597 11069 12631
rect 11103 12628 11115 12631
rect 12342 12628 12348 12640
rect 11103 12600 12348 12628
rect 11103 12597 11115 12600
rect 11057 12591 11115 12597
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 13357 12631 13415 12637
rect 13357 12628 13369 12631
rect 12584 12600 13369 12628
rect 12584 12588 12590 12600
rect 13357 12597 13369 12600
rect 13403 12597 13415 12631
rect 13357 12591 13415 12597
rect 15105 12631 15163 12637
rect 15105 12597 15117 12631
rect 15151 12628 15163 12631
rect 15470 12628 15476 12640
rect 15151 12600 15476 12628
rect 15151 12597 15163 12600
rect 15105 12591 15163 12597
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 15580 12628 15608 12668
rect 16040 12668 16313 12696
rect 16040 12628 16068 12668
rect 16301 12665 16313 12668
rect 16347 12665 16359 12699
rect 16301 12659 16359 12665
rect 22370 12656 22376 12708
rect 22428 12656 22434 12708
rect 24210 12656 24216 12708
rect 24268 12696 24274 12708
rect 29840 12696 29868 12736
rect 31754 12724 31760 12736
rect 31812 12724 31818 12776
rect 24268 12668 29868 12696
rect 31864 12696 31892 12804
rect 32769 12801 32781 12835
rect 32815 12801 32827 12835
rect 32769 12795 32827 12801
rect 32784 12764 32812 12795
rect 33042 12792 33048 12844
rect 33100 12792 33106 12844
rect 33152 12841 33180 12872
rect 34885 12869 34897 12903
rect 34931 12900 34943 12903
rect 35618 12900 35624 12912
rect 34931 12872 35624 12900
rect 34931 12869 34943 12872
rect 34885 12863 34943 12869
rect 35618 12860 35624 12872
rect 35676 12860 35682 12912
rect 33137 12835 33195 12841
rect 33137 12801 33149 12835
rect 33183 12801 33195 12835
rect 33137 12795 33195 12801
rect 33318 12792 33324 12844
rect 33376 12832 33382 12844
rect 33781 12835 33839 12841
rect 33781 12832 33793 12835
rect 33376 12804 33793 12832
rect 33376 12792 33382 12804
rect 33781 12801 33793 12804
rect 33827 12832 33839 12835
rect 33962 12832 33968 12844
rect 33827 12804 33968 12832
rect 33827 12801 33839 12804
rect 33781 12795 33839 12801
rect 33962 12792 33968 12804
rect 34020 12792 34026 12844
rect 34793 12835 34851 12841
rect 34793 12801 34805 12835
rect 34839 12801 34851 12835
rect 34793 12795 34851 12801
rect 32858 12764 32864 12776
rect 32784 12736 32864 12764
rect 32858 12724 32864 12736
rect 32916 12764 32922 12776
rect 34808 12764 34836 12795
rect 35250 12792 35256 12844
rect 35308 12832 35314 12844
rect 35713 12835 35771 12841
rect 35713 12832 35725 12835
rect 35308 12804 35725 12832
rect 35308 12792 35314 12804
rect 35713 12801 35725 12804
rect 35759 12801 35771 12835
rect 35713 12795 35771 12801
rect 37458 12792 37464 12844
rect 37516 12832 37522 12844
rect 37553 12835 37611 12841
rect 37553 12832 37565 12835
rect 37516 12804 37565 12832
rect 37516 12792 37522 12804
rect 37553 12801 37565 12804
rect 37599 12801 37611 12835
rect 37553 12795 37611 12801
rect 37826 12792 37832 12844
rect 37884 12832 37890 12844
rect 38197 12835 38255 12841
rect 38197 12832 38209 12835
rect 37884 12804 38209 12832
rect 37884 12792 37890 12804
rect 38197 12801 38209 12804
rect 38243 12801 38255 12835
rect 38197 12795 38255 12801
rect 32916 12736 34836 12764
rect 32916 12724 32922 12736
rect 34882 12724 34888 12776
rect 34940 12764 34946 12776
rect 34977 12767 35035 12773
rect 34977 12764 34989 12767
rect 34940 12736 34989 12764
rect 34940 12724 34946 12736
rect 34977 12733 34989 12736
rect 35023 12764 35035 12767
rect 35989 12767 36047 12773
rect 35989 12764 36001 12767
rect 35023 12736 36001 12764
rect 35023 12733 35035 12736
rect 34977 12727 35035 12733
rect 35989 12733 36001 12736
rect 36035 12733 36047 12767
rect 35989 12727 36047 12733
rect 37645 12699 37703 12705
rect 37645 12696 37657 12699
rect 31864 12668 37657 12696
rect 24268 12656 24274 12668
rect 37645 12665 37657 12668
rect 37691 12665 37703 12699
rect 37645 12659 37703 12665
rect 15580 12600 16068 12628
rect 16117 12631 16175 12637
rect 16117 12597 16129 12631
rect 16163 12628 16175 12631
rect 16574 12628 16580 12640
rect 16163 12600 16580 12628
rect 16163 12597 16175 12600
rect 16117 12591 16175 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 16942 12588 16948 12640
rect 17000 12628 17006 12640
rect 17770 12628 17776 12640
rect 17000 12600 17776 12628
rect 17000 12588 17006 12600
rect 17770 12588 17776 12600
rect 17828 12588 17834 12640
rect 18322 12588 18328 12640
rect 18380 12628 18386 12640
rect 18598 12628 18604 12640
rect 18380 12600 18604 12628
rect 18380 12588 18386 12600
rect 18598 12588 18604 12600
rect 18656 12588 18662 12640
rect 20438 12588 20444 12640
rect 20496 12628 20502 12640
rect 24673 12631 24731 12637
rect 24673 12628 24685 12631
rect 20496 12600 24685 12628
rect 20496 12588 20502 12600
rect 24673 12597 24685 12600
rect 24719 12597 24731 12631
rect 24673 12591 24731 12597
rect 25498 12588 25504 12640
rect 25556 12628 25562 12640
rect 25682 12628 25688 12640
rect 25556 12600 25688 12628
rect 25556 12588 25562 12600
rect 25682 12588 25688 12600
rect 25740 12588 25746 12640
rect 25866 12588 25872 12640
rect 25924 12628 25930 12640
rect 27430 12628 27436 12640
rect 25924 12600 27436 12628
rect 25924 12588 25930 12600
rect 27430 12588 27436 12600
rect 27488 12588 27494 12640
rect 29273 12631 29331 12637
rect 29273 12597 29285 12631
rect 29319 12628 29331 12631
rect 30742 12628 30748 12640
rect 29319 12600 30748 12628
rect 29319 12597 29331 12600
rect 29273 12591 29331 12597
rect 30742 12588 30748 12600
rect 30800 12588 30806 12640
rect 33318 12588 33324 12640
rect 33376 12588 33382 12640
rect 33870 12588 33876 12640
rect 33928 12588 33934 12640
rect 34146 12588 34152 12640
rect 34204 12628 34210 12640
rect 34425 12631 34483 12637
rect 34425 12628 34437 12631
rect 34204 12600 34437 12628
rect 34204 12588 34210 12600
rect 34425 12597 34437 12600
rect 34471 12597 34483 12631
rect 34425 12591 34483 12597
rect 34882 12588 34888 12640
rect 34940 12628 34946 12640
rect 35250 12628 35256 12640
rect 34940 12600 35256 12628
rect 34940 12588 34946 12600
rect 35250 12588 35256 12600
rect 35308 12588 35314 12640
rect 38286 12588 38292 12640
rect 38344 12588 38350 12640
rect 1104 12538 39192 12560
rect 1104 12486 5711 12538
rect 5763 12486 5775 12538
rect 5827 12486 5839 12538
rect 5891 12486 5903 12538
rect 5955 12486 5967 12538
rect 6019 12486 15233 12538
rect 15285 12486 15297 12538
rect 15349 12486 15361 12538
rect 15413 12486 15425 12538
rect 15477 12486 15489 12538
rect 15541 12486 24755 12538
rect 24807 12486 24819 12538
rect 24871 12486 24883 12538
rect 24935 12486 24947 12538
rect 24999 12486 25011 12538
rect 25063 12486 34277 12538
rect 34329 12486 34341 12538
rect 34393 12486 34405 12538
rect 34457 12486 34469 12538
rect 34521 12486 34533 12538
rect 34585 12486 39192 12538
rect 1104 12464 39192 12486
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 3602 12424 3608 12436
rect 1820 12396 3608 12424
rect 1820 12384 1826 12396
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 9950 12424 9956 12436
rect 4080 12396 9956 12424
rect 4080 12356 4108 12396
rect 9950 12384 9956 12396
rect 10008 12424 10014 12436
rect 10226 12424 10232 12436
rect 10008 12396 10232 12424
rect 10008 12384 10014 12396
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 10594 12384 10600 12436
rect 10652 12424 10658 12436
rect 10652 12396 12434 12424
rect 10652 12384 10658 12396
rect 1964 12328 4108 12356
rect 5721 12359 5779 12365
rect 1964 12229 1992 12328
rect 5721 12325 5733 12359
rect 5767 12356 5779 12359
rect 5767 12328 7696 12356
rect 5767 12325 5779 12328
rect 5721 12319 5779 12325
rect 2038 12248 2044 12300
rect 2096 12248 2102 12300
rect 3142 12248 3148 12300
rect 3200 12288 3206 12300
rect 5736 12288 5764 12319
rect 3200 12260 5764 12288
rect 3200 12248 3206 12260
rect 5810 12248 5816 12300
rect 5868 12288 5874 12300
rect 7006 12288 7012 12300
rect 5868 12260 7012 12288
rect 5868 12248 5874 12260
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12288 7527 12291
rect 7668 12288 7696 12328
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 9122 12356 9128 12368
rect 8996 12328 9128 12356
rect 8996 12316 9002 12328
rect 9122 12316 9128 12328
rect 9180 12316 9186 12368
rect 9769 12359 9827 12365
rect 9769 12325 9781 12359
rect 9815 12356 9827 12359
rect 10778 12356 10784 12368
rect 9815 12328 10784 12356
rect 9815 12325 9827 12328
rect 9769 12319 9827 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 11057 12359 11115 12365
rect 11057 12325 11069 12359
rect 11103 12356 11115 12359
rect 11238 12356 11244 12368
rect 11103 12328 11244 12356
rect 11103 12325 11115 12328
rect 11057 12319 11115 12325
rect 11238 12316 11244 12328
rect 11296 12316 11302 12368
rect 12406 12356 12434 12396
rect 12526 12384 12532 12436
rect 12584 12384 12590 12436
rect 13722 12384 13728 12436
rect 13780 12384 13786 12436
rect 15473 12427 15531 12433
rect 15473 12393 15485 12427
rect 15519 12424 15531 12427
rect 15562 12424 15568 12436
rect 15519 12396 15568 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 16025 12427 16083 12433
rect 16025 12393 16037 12427
rect 16071 12424 16083 12427
rect 16390 12424 16396 12436
rect 16071 12396 16396 12424
rect 16071 12393 16083 12396
rect 16025 12387 16083 12393
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16500 12396 16712 12424
rect 12713 12359 12771 12365
rect 12713 12356 12725 12359
rect 12406 12328 12725 12356
rect 12713 12325 12725 12328
rect 12759 12325 12771 12359
rect 16500 12356 16528 12396
rect 12713 12319 12771 12325
rect 13188 12328 16528 12356
rect 16684 12356 16712 12396
rect 17770 12384 17776 12436
rect 17828 12384 17834 12436
rect 20346 12384 20352 12436
rect 20404 12384 20410 12436
rect 21082 12384 21088 12436
rect 21140 12384 21146 12436
rect 21266 12384 21272 12436
rect 21324 12384 21330 12436
rect 23106 12424 23112 12436
rect 21376 12396 23112 12424
rect 17218 12356 17224 12368
rect 16684 12328 17224 12356
rect 7515 12260 7604 12288
rect 7668 12260 12388 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12189 2007 12223
rect 2056 12220 2084 12248
rect 2590 12220 2596 12232
rect 2056 12192 2596 12220
rect 1949 12183 2007 12189
rect 2590 12180 2596 12192
rect 2648 12220 2654 12232
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 2648 12192 3249 12220
rect 2648 12180 2654 12192
rect 3237 12189 3249 12192
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 3970 12180 3976 12232
rect 4028 12180 4034 12232
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 5684 12192 6285 12220
rect 5684 12180 5690 12192
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 2041 12155 2099 12161
rect 2041 12121 2053 12155
rect 2087 12152 2099 12155
rect 2087 12124 3740 12152
rect 2087 12121 2099 12124
rect 2041 12115 2099 12121
rect 2682 12044 2688 12096
rect 2740 12044 2746 12096
rect 3234 12044 3240 12096
rect 3292 12084 3298 12096
rect 3329 12087 3387 12093
rect 3329 12084 3341 12087
rect 3292 12056 3341 12084
rect 3292 12044 3298 12056
rect 3329 12053 3341 12056
rect 3375 12053 3387 12087
rect 3712 12084 3740 12124
rect 3878 12112 3884 12164
rect 3936 12152 3942 12164
rect 4249 12155 4307 12161
rect 4249 12152 4261 12155
rect 3936 12124 4261 12152
rect 3936 12112 3942 12124
rect 4249 12121 4261 12124
rect 4295 12121 4307 12155
rect 4249 12115 4307 12121
rect 4356 12124 4738 12152
rect 4356 12084 4384 12124
rect 7374 12112 7380 12164
rect 7432 12112 7438 12164
rect 7576 12152 7604 12260
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 7800 12192 8401 12220
rect 7800 12180 7806 12192
rect 8389 12189 8401 12192
rect 8435 12220 8447 12223
rect 8938 12220 8944 12232
rect 8435 12192 8944 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8938 12180 8944 12192
rect 8996 12220 9002 12232
rect 9677 12223 9735 12229
rect 8996 12192 9536 12220
rect 8996 12180 9002 12192
rect 7834 12152 7840 12164
rect 7576 12124 7840 12152
rect 7834 12112 7840 12124
rect 7892 12112 7898 12164
rect 9398 12152 9404 12164
rect 8404 12124 9404 12152
rect 3712 12056 4384 12084
rect 3329 12047 3387 12053
rect 6178 12044 6184 12096
rect 6236 12084 6242 12096
rect 6365 12087 6423 12093
rect 6365 12084 6377 12087
rect 6236 12056 6377 12084
rect 6236 12044 6242 12056
rect 6365 12053 6377 12056
rect 6411 12053 6423 12087
rect 6365 12047 6423 12053
rect 6454 12044 6460 12096
rect 6512 12084 6518 12096
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6512 12056 6929 12084
rect 6512 12044 6518 12056
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 6917 12047 6975 12053
rect 7285 12087 7343 12093
rect 7285 12053 7297 12087
rect 7331 12084 7343 12087
rect 8404 12084 8432 12124
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 9508 12152 9536 12192
rect 9677 12189 9689 12223
rect 9723 12220 9735 12223
rect 9858 12220 9864 12232
rect 9723 12192 9864 12220
rect 9723 12189 9735 12192
rect 9677 12183 9735 12189
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10502 12220 10508 12232
rect 10367 12192 10508 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10502 12180 10508 12192
rect 10560 12220 10566 12232
rect 11238 12220 11244 12232
rect 10560 12192 11244 12220
rect 10560 12180 10566 12192
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 11480 12192 11529 12220
rect 11480 12180 11486 12192
rect 11517 12189 11529 12192
rect 11563 12220 11575 12223
rect 11882 12220 11888 12232
rect 11563 12192 11888 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 9950 12152 9956 12164
rect 9508 12124 9956 12152
rect 9950 12112 9956 12124
rect 10008 12112 10014 12164
rect 10594 12152 10600 12164
rect 10060 12124 10600 12152
rect 7331 12056 8432 12084
rect 8481 12087 8539 12093
rect 7331 12053 7343 12056
rect 7285 12047 7343 12053
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 8662 12084 8668 12096
rect 8527 12056 8668 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10060 12084 10088 12124
rect 10594 12112 10600 12124
rect 10652 12112 10658 12164
rect 12360 12161 12388 12260
rect 13188 12229 13216 12328
rect 17218 12316 17224 12328
rect 17276 12316 17282 12368
rect 17310 12316 17316 12368
rect 17368 12356 17374 12368
rect 17368 12328 17540 12356
rect 17368 12316 17374 12328
rect 13372 12260 16436 12288
rect 13372 12232 13400 12260
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 13354 12180 13360 12232
rect 13412 12180 13418 12232
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 14056 12192 14289 12220
rect 14056 12180 14062 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 14734 12180 14740 12232
rect 14792 12180 14798 12232
rect 14826 12180 14832 12232
rect 14884 12220 14890 12232
rect 14921 12223 14979 12229
rect 14921 12220 14933 12223
rect 14884 12192 14933 12220
rect 14884 12180 14890 12192
rect 14921 12189 14933 12192
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 15286 12180 15292 12232
rect 15344 12180 15350 12232
rect 16408 12220 16436 12260
rect 16482 12248 16488 12300
rect 16540 12248 16546 12300
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12288 16727 12291
rect 16758 12288 16764 12300
rect 16715 12260 16764 12288
rect 16715 12257 16727 12260
rect 16669 12251 16727 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 17402 12288 17408 12300
rect 17236 12260 17408 12288
rect 17236 12229 17264 12260
rect 17402 12248 17408 12260
rect 17460 12248 17466 12300
rect 17512 12229 17540 12328
rect 17678 12316 17684 12368
rect 17736 12356 17742 12368
rect 17954 12356 17960 12368
rect 17736 12328 17960 12356
rect 17736 12316 17742 12328
rect 17954 12316 17960 12328
rect 18012 12316 18018 12368
rect 19702 12356 19708 12368
rect 18616 12328 19708 12356
rect 18616 12297 18644 12328
rect 19702 12316 19708 12328
rect 19760 12316 19766 12368
rect 20238 12359 20296 12365
rect 20238 12325 20250 12359
rect 20284 12356 20296 12359
rect 21100 12356 21128 12384
rect 20284 12328 21128 12356
rect 20284 12325 20296 12328
rect 20238 12319 20296 12325
rect 18601 12291 18659 12297
rect 18601 12257 18613 12291
rect 18647 12257 18659 12291
rect 18601 12251 18659 12257
rect 18690 12248 18696 12300
rect 18748 12248 18754 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 20441 12291 20499 12297
rect 20441 12288 20453 12291
rect 19392 12260 20453 12288
rect 19392 12248 19398 12260
rect 20441 12257 20453 12260
rect 20487 12257 20499 12291
rect 20441 12251 20499 12257
rect 20809 12291 20867 12297
rect 20809 12257 20821 12291
rect 20855 12288 20867 12291
rect 21376 12288 21404 12396
rect 23106 12384 23112 12396
rect 23164 12384 23170 12436
rect 23658 12384 23664 12436
rect 23716 12424 23722 12436
rect 26050 12424 26056 12436
rect 23716 12396 26056 12424
rect 23716 12384 23722 12396
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 26694 12384 26700 12436
rect 26752 12424 26758 12436
rect 27430 12424 27436 12436
rect 26752 12396 27436 12424
rect 26752 12384 26758 12396
rect 27430 12384 27436 12396
rect 27488 12424 27494 12436
rect 28994 12424 29000 12436
rect 27488 12396 29000 12424
rect 27488 12384 27494 12396
rect 21450 12316 21456 12368
rect 21508 12356 21514 12368
rect 21634 12356 21640 12368
rect 21508 12328 21640 12356
rect 21508 12316 21514 12328
rect 21634 12316 21640 12328
rect 21692 12316 21698 12368
rect 21821 12291 21879 12297
rect 21821 12288 21833 12291
rect 20855 12260 21404 12288
rect 21468 12260 21833 12288
rect 20855 12257 20867 12260
rect 20809 12251 20867 12257
rect 17221 12223 17279 12229
rect 16408 12214 16620 12220
rect 16408 12192 16712 12214
rect 16592 12186 16712 12192
rect 11057 12155 11115 12161
rect 11057 12121 11069 12155
rect 11103 12152 11115 12155
rect 12345 12155 12403 12161
rect 11103 12124 11928 12152
rect 11103 12121 11115 12124
rect 11057 12115 11115 12121
rect 9732 12056 10088 12084
rect 9732 12044 9738 12056
rect 10226 12044 10232 12096
rect 10284 12084 10290 12096
rect 10413 12087 10471 12093
rect 10413 12084 10425 12087
rect 10284 12056 10425 12084
rect 10284 12044 10290 12056
rect 10413 12053 10425 12056
rect 10459 12053 10471 12087
rect 10413 12047 10471 12053
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 11146 12084 11152 12096
rect 10836 12056 11152 12084
rect 10836 12044 10842 12056
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 11606 12044 11612 12096
rect 11664 12044 11670 12096
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 11793 12087 11851 12093
rect 11793 12084 11805 12087
rect 11756 12056 11805 12084
rect 11756 12044 11762 12056
rect 11793 12053 11805 12056
rect 11839 12053 11851 12087
rect 11900 12084 11928 12124
rect 12345 12121 12357 12155
rect 12391 12121 12403 12155
rect 12345 12115 12403 12121
rect 12561 12155 12619 12161
rect 12561 12121 12573 12155
rect 12607 12152 12619 12155
rect 13262 12152 13268 12164
rect 12607 12124 13268 12152
rect 12607 12121 12619 12124
rect 12561 12115 12619 12121
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 13449 12155 13507 12161
rect 13449 12121 13461 12155
rect 13495 12152 13507 12155
rect 13630 12152 13636 12164
rect 13495 12124 13636 12152
rect 13495 12121 13507 12124
rect 13449 12115 13507 12121
rect 13630 12112 13636 12124
rect 13688 12112 13694 12164
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 14752 12152 14780 12180
rect 15105 12155 15163 12161
rect 15105 12152 15117 12155
rect 13780 12124 15117 12152
rect 13780 12112 13786 12124
rect 15105 12121 15117 12124
rect 15151 12121 15163 12155
rect 15105 12115 15163 12121
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12152 15255 12155
rect 16206 12152 16212 12164
rect 15243 12124 16212 12152
rect 15243 12121 15255 12124
rect 15197 12115 15255 12121
rect 16206 12112 16212 12124
rect 16264 12112 16270 12164
rect 16684 12152 16712 12186
rect 17221 12189 17233 12223
rect 17267 12189 17279 12223
rect 17221 12183 17279 12189
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12220 17647 12223
rect 17678 12220 17684 12232
rect 17635 12192 17684 12220
rect 17635 12189 17647 12192
rect 17589 12183 17647 12189
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12220 18475 12223
rect 18708 12220 18736 12248
rect 18463 12192 18736 12220
rect 19429 12223 19487 12229
rect 18463 12189 18475 12192
rect 18417 12183 18475 12189
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12220 20131 12223
rect 20530 12220 20536 12232
rect 20119 12192 20536 12220
rect 20119 12189 20131 12192
rect 20073 12183 20131 12189
rect 17405 12155 17463 12161
rect 17405 12152 17417 12155
rect 16684 12124 17417 12152
rect 17405 12121 17417 12124
rect 17451 12152 17463 12155
rect 17862 12152 17868 12164
rect 17451 12124 17868 12152
rect 17451 12121 17463 12124
rect 17405 12115 17463 12121
rect 17862 12112 17868 12124
rect 17920 12112 17926 12164
rect 13906 12084 13912 12096
rect 11900 12056 13912 12084
rect 11793 12047 11851 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14369 12087 14427 12093
rect 14369 12053 14381 12087
rect 14415 12084 14427 12087
rect 14734 12084 14740 12096
rect 14415 12056 14740 12084
rect 14415 12053 14427 12056
rect 14369 12047 14427 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16393 12087 16451 12093
rect 16393 12084 16405 12087
rect 16080 12056 16405 12084
rect 16080 12044 16086 12056
rect 16393 12053 16405 12056
rect 16439 12053 16451 12087
rect 16393 12047 16451 12053
rect 16758 12044 16764 12096
rect 16816 12084 16822 12096
rect 18414 12084 18420 12096
rect 16816 12056 18420 12084
rect 16816 12044 16822 12056
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 19444 12084 19472 12183
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 21468 12220 21496 12260
rect 21821 12257 21833 12260
rect 21867 12257 21879 12291
rect 21821 12251 21879 12257
rect 25130 12248 25136 12300
rect 25188 12288 25194 12300
rect 25685 12291 25743 12297
rect 25685 12288 25697 12291
rect 25188 12260 25697 12288
rect 25188 12248 25194 12260
rect 25685 12257 25697 12260
rect 25731 12288 25743 12291
rect 25958 12288 25964 12300
rect 25731 12260 25964 12288
rect 25731 12257 25743 12260
rect 25685 12251 25743 12257
rect 25958 12248 25964 12260
rect 26016 12248 26022 12300
rect 20772 12192 21496 12220
rect 20772 12180 20778 12192
rect 21634 12180 21640 12232
rect 21692 12220 21698 12232
rect 22465 12223 22523 12229
rect 22465 12220 22477 12223
rect 21692 12192 22477 12220
rect 21692 12180 21698 12192
rect 22465 12189 22477 12192
rect 22511 12189 22523 12223
rect 22465 12183 22523 12189
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 23198 12220 23204 12232
rect 22704 12192 23204 12220
rect 22704 12180 22710 12192
rect 23198 12180 23204 12192
rect 23256 12180 23262 12232
rect 23842 12180 23848 12232
rect 23900 12220 23906 12232
rect 24486 12220 24492 12232
rect 23900 12192 24492 12220
rect 23900 12180 23906 12192
rect 24486 12180 24492 12192
rect 24544 12180 24550 12232
rect 24578 12180 24584 12232
rect 24636 12220 24642 12232
rect 24857 12223 24915 12229
rect 24857 12220 24869 12223
rect 24636 12192 24869 12220
rect 24636 12180 24642 12192
rect 24857 12189 24869 12192
rect 24903 12189 24915 12223
rect 24857 12183 24915 12189
rect 27338 12180 27344 12232
rect 27396 12220 27402 12232
rect 27890 12220 27896 12232
rect 27396 12192 27896 12220
rect 27396 12180 27402 12192
rect 27890 12180 27896 12192
rect 27948 12180 27954 12232
rect 28276 12229 28304 12396
rect 28994 12384 29000 12396
rect 29052 12384 29058 12436
rect 31110 12384 31116 12436
rect 31168 12424 31174 12436
rect 32585 12427 32643 12433
rect 32585 12424 32597 12427
rect 31168 12396 32597 12424
rect 31168 12384 31174 12396
rect 32585 12393 32597 12396
rect 32631 12393 32643 12427
rect 32585 12387 32643 12393
rect 33042 12384 33048 12436
rect 33100 12424 33106 12436
rect 34882 12424 34888 12436
rect 33100 12396 34888 12424
rect 33100 12384 33106 12396
rect 34882 12384 34888 12396
rect 34940 12384 34946 12436
rect 35066 12384 35072 12436
rect 35124 12384 35130 12436
rect 35986 12384 35992 12436
rect 36044 12384 36050 12436
rect 37182 12384 37188 12436
rect 37240 12424 37246 12436
rect 37921 12427 37979 12433
rect 37921 12424 37933 12427
rect 37240 12396 37933 12424
rect 37240 12384 37246 12396
rect 37921 12393 37933 12396
rect 37967 12393 37979 12427
rect 37921 12387 37979 12393
rect 31662 12316 31668 12368
rect 31720 12356 31726 12368
rect 32769 12359 32827 12365
rect 32769 12356 32781 12359
rect 31720 12328 32781 12356
rect 31720 12316 31726 12328
rect 32769 12325 32781 12328
rect 32815 12325 32827 12359
rect 32769 12319 32827 12325
rect 33134 12316 33140 12368
rect 33192 12356 33198 12368
rect 36817 12359 36875 12365
rect 36817 12356 36829 12359
rect 33192 12328 36829 12356
rect 33192 12316 33198 12328
rect 36817 12325 36829 12328
rect 36863 12325 36875 12359
rect 36817 12319 36875 12325
rect 28350 12248 28356 12300
rect 28408 12288 28414 12300
rect 28537 12291 28595 12297
rect 28537 12288 28549 12291
rect 28408 12260 28549 12288
rect 28408 12248 28414 12260
rect 28537 12257 28549 12260
rect 28583 12288 28595 12291
rect 28626 12288 28632 12300
rect 28583 12260 28632 12288
rect 28583 12257 28595 12260
rect 28537 12251 28595 12257
rect 28626 12248 28632 12260
rect 28684 12248 28690 12300
rect 29362 12248 29368 12300
rect 29420 12288 29426 12300
rect 30193 12291 30251 12297
rect 30193 12288 30205 12291
rect 29420 12260 30205 12288
rect 29420 12248 29426 12260
rect 30193 12257 30205 12260
rect 30239 12257 30251 12291
rect 30193 12251 30251 12257
rect 30469 12291 30527 12297
rect 30469 12257 30481 12291
rect 30515 12288 30527 12291
rect 31754 12288 31760 12300
rect 30515 12260 31760 12288
rect 30515 12257 30527 12260
rect 30469 12251 30527 12257
rect 31754 12248 31760 12260
rect 31812 12248 31818 12300
rect 31941 12291 31999 12297
rect 31941 12257 31953 12291
rect 31987 12288 31999 12291
rect 32858 12288 32864 12300
rect 31987 12260 32864 12288
rect 31987 12257 31999 12260
rect 31941 12251 31999 12257
rect 32858 12248 32864 12260
rect 32916 12248 32922 12300
rect 33410 12248 33416 12300
rect 33468 12288 33474 12300
rect 33686 12288 33692 12300
rect 33468 12260 33692 12288
rect 33468 12248 33474 12260
rect 33686 12248 33692 12260
rect 33744 12288 33750 12300
rect 33781 12291 33839 12297
rect 33781 12288 33793 12291
rect 33744 12260 33793 12288
rect 33744 12248 33750 12260
rect 33781 12257 33793 12260
rect 33827 12257 33839 12291
rect 33781 12251 33839 12257
rect 35066 12248 35072 12300
rect 35124 12288 35130 12300
rect 37458 12288 37464 12300
rect 35124 12260 37464 12288
rect 35124 12248 35130 12260
rect 28261 12223 28319 12229
rect 28261 12189 28273 12223
rect 28307 12189 28319 12223
rect 31602 12192 34560 12220
rect 28261 12183 28319 12189
rect 19521 12155 19579 12161
rect 19521 12121 19533 12155
rect 19567 12152 19579 12155
rect 20806 12152 20812 12164
rect 19567 12124 20812 12152
rect 19567 12121 19579 12124
rect 19521 12115 19579 12121
rect 20806 12112 20812 12124
rect 20864 12112 20870 12164
rect 20990 12112 20996 12164
rect 21048 12152 21054 12164
rect 21542 12152 21548 12164
rect 21048 12124 21548 12152
rect 21048 12112 21054 12124
rect 21542 12112 21548 12124
rect 21600 12152 21606 12164
rect 21729 12155 21787 12161
rect 21729 12152 21741 12155
rect 21600 12124 21741 12152
rect 21600 12112 21606 12124
rect 21729 12121 21741 12124
rect 21775 12121 21787 12155
rect 21729 12115 21787 12121
rect 22554 12112 22560 12164
rect 22612 12152 22618 12164
rect 22741 12155 22799 12161
rect 22741 12152 22753 12155
rect 22612 12124 22753 12152
rect 22612 12112 22618 12124
rect 22741 12121 22753 12124
rect 22787 12121 22799 12155
rect 22741 12115 22799 12121
rect 23014 12112 23020 12164
rect 23072 12152 23078 12164
rect 25406 12152 25412 12164
rect 23072 12124 25412 12152
rect 23072 12112 23078 12124
rect 24504 12096 24532 12124
rect 25406 12112 25412 12124
rect 25464 12112 25470 12164
rect 25961 12155 26019 12161
rect 25961 12121 25973 12155
rect 26007 12121 26019 12155
rect 27246 12152 27252 12164
rect 27186 12124 27252 12152
rect 25961 12115 26019 12121
rect 20622 12084 20628 12096
rect 19444 12056 20628 12084
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 21082 12044 21088 12096
rect 21140 12084 21146 12096
rect 21450 12084 21456 12096
rect 21140 12056 21456 12084
rect 21140 12044 21146 12056
rect 21450 12044 21456 12056
rect 21508 12084 21514 12096
rect 21637 12087 21695 12093
rect 21637 12084 21649 12087
rect 21508 12056 21649 12084
rect 21508 12044 21514 12056
rect 21637 12053 21649 12056
rect 21683 12053 21695 12087
rect 21637 12047 21695 12053
rect 21818 12044 21824 12096
rect 21876 12084 21882 12096
rect 23937 12087 23995 12093
rect 23937 12084 23949 12087
rect 21876 12056 23949 12084
rect 21876 12044 21882 12056
rect 23937 12053 23949 12056
rect 23983 12053 23995 12087
rect 23937 12047 23995 12053
rect 24486 12044 24492 12096
rect 24544 12044 24550 12096
rect 24949 12087 25007 12093
rect 24949 12053 24961 12087
rect 24995 12084 25007 12087
rect 25682 12084 25688 12096
rect 24995 12056 25688 12084
rect 24995 12053 25007 12056
rect 24949 12047 25007 12053
rect 25682 12044 25688 12056
rect 25740 12044 25746 12096
rect 25976 12084 26004 12115
rect 27246 12112 27252 12124
rect 27304 12112 27310 12164
rect 29270 12112 29276 12164
rect 29328 12152 29334 12164
rect 30006 12152 30012 12164
rect 29328 12124 30012 12152
rect 29328 12112 29334 12124
rect 30006 12112 30012 12124
rect 30064 12112 30070 12164
rect 32401 12155 32459 12161
rect 32401 12152 32413 12155
rect 31864 12124 32413 12152
rect 26970 12084 26976 12096
rect 25976 12056 26976 12084
rect 26970 12044 26976 12056
rect 27028 12044 27034 12096
rect 27338 12044 27344 12096
rect 27396 12084 27402 12096
rect 27433 12087 27491 12093
rect 27433 12084 27445 12087
rect 27396 12056 27445 12084
rect 27396 12044 27402 12056
rect 27433 12053 27445 12056
rect 27479 12053 27491 12087
rect 27433 12047 27491 12053
rect 27522 12044 27528 12096
rect 27580 12084 27586 12096
rect 27893 12087 27951 12093
rect 27893 12084 27905 12087
rect 27580 12056 27905 12084
rect 27580 12044 27586 12056
rect 27893 12053 27905 12056
rect 27939 12053 27951 12087
rect 27893 12047 27951 12053
rect 28353 12087 28411 12093
rect 28353 12053 28365 12087
rect 28399 12084 28411 12087
rect 28718 12084 28724 12096
rect 28399 12056 28724 12084
rect 28399 12053 28411 12056
rect 28353 12047 28411 12053
rect 28718 12044 28724 12056
rect 28776 12084 28782 12096
rect 28902 12084 28908 12096
rect 28776 12056 28908 12084
rect 28776 12044 28782 12056
rect 28902 12044 28908 12056
rect 28960 12044 28966 12096
rect 29914 12044 29920 12096
rect 29972 12084 29978 12096
rect 30374 12084 30380 12096
rect 29972 12056 30380 12084
rect 29972 12044 29978 12056
rect 30374 12044 30380 12056
rect 30432 12044 30438 12096
rect 30558 12044 30564 12096
rect 30616 12084 30622 12096
rect 31386 12084 31392 12096
rect 30616 12056 31392 12084
rect 30616 12044 30622 12056
rect 31386 12044 31392 12056
rect 31444 12044 31450 12096
rect 31478 12044 31484 12096
rect 31536 12084 31542 12096
rect 31864 12084 31892 12124
rect 32401 12121 32413 12124
rect 32447 12121 32459 12155
rect 32766 12152 32772 12164
rect 32401 12115 32459 12121
rect 32508 12124 32772 12152
rect 31536 12056 31892 12084
rect 31536 12044 31542 12056
rect 32306 12044 32312 12096
rect 32364 12084 32370 12096
rect 32508 12084 32536 12124
rect 32766 12112 32772 12124
rect 32824 12152 32830 12164
rect 33042 12152 33048 12164
rect 32824 12124 33048 12152
rect 32824 12112 32830 12124
rect 33042 12112 33048 12124
rect 33100 12112 33106 12164
rect 33134 12112 33140 12164
rect 33192 12152 33198 12164
rect 33597 12155 33655 12161
rect 33597 12152 33609 12155
rect 33192 12124 33609 12152
rect 33192 12112 33198 12124
rect 33597 12121 33609 12124
rect 33643 12121 33655 12155
rect 33597 12115 33655 12121
rect 33689 12155 33747 12161
rect 33689 12121 33701 12155
rect 33735 12152 33747 12155
rect 34146 12152 34152 12164
rect 33735 12124 34152 12152
rect 33735 12121 33747 12124
rect 33689 12115 33747 12121
rect 34146 12112 34152 12124
rect 34204 12112 34210 12164
rect 32364 12056 32536 12084
rect 32364 12044 32370 12056
rect 32582 12044 32588 12096
rect 32640 12093 32646 12096
rect 32640 12087 32659 12093
rect 32647 12053 32659 12087
rect 32640 12047 32659 12053
rect 32640 12044 32646 12047
rect 32858 12044 32864 12096
rect 32916 12084 32922 12096
rect 33229 12087 33287 12093
rect 33229 12084 33241 12087
rect 32916 12056 33241 12084
rect 32916 12044 32922 12056
rect 33229 12053 33241 12056
rect 33275 12053 33287 12087
rect 34532 12084 34560 12192
rect 34606 12180 34612 12232
rect 34664 12220 34670 12232
rect 35805 12223 35863 12229
rect 35805 12220 35817 12223
rect 34664 12192 35817 12220
rect 34664 12180 34670 12192
rect 35805 12189 35817 12192
rect 35851 12189 35863 12223
rect 35805 12183 35863 12189
rect 35894 12180 35900 12232
rect 35952 12180 35958 12232
rect 36740 12229 36768 12260
rect 37458 12248 37464 12260
rect 37516 12248 37522 12300
rect 36725 12223 36783 12229
rect 36725 12189 36737 12223
rect 36771 12189 36783 12223
rect 37476 12220 37504 12248
rect 37829 12223 37887 12229
rect 37829 12220 37841 12223
rect 37476 12192 37841 12220
rect 36725 12183 36783 12189
rect 37829 12189 37841 12192
rect 37875 12220 37887 12223
rect 38010 12220 38016 12232
rect 37875 12192 38016 12220
rect 37875 12189 37887 12192
rect 37829 12183 37887 12189
rect 38010 12180 38016 12192
rect 38068 12180 38074 12232
rect 38378 12180 38384 12232
rect 38436 12220 38442 12232
rect 38473 12223 38531 12229
rect 38473 12220 38485 12223
rect 38436 12192 38485 12220
rect 38436 12180 38442 12192
rect 38473 12189 38485 12192
rect 38519 12189 38531 12223
rect 38473 12183 38531 12189
rect 34790 12112 34796 12164
rect 34848 12152 34854 12164
rect 34977 12155 35035 12161
rect 34977 12152 34989 12155
rect 34848 12124 34989 12152
rect 34848 12112 34854 12124
rect 34977 12121 34989 12124
rect 35023 12121 35035 12155
rect 34977 12115 35035 12121
rect 35158 12112 35164 12164
rect 35216 12152 35222 12164
rect 38565 12155 38623 12161
rect 38565 12152 38577 12155
rect 35216 12124 38577 12152
rect 35216 12112 35222 12124
rect 38565 12121 38577 12124
rect 38611 12121 38623 12155
rect 38565 12115 38623 12121
rect 36078 12084 36084 12096
rect 34532 12056 36084 12084
rect 33229 12047 33287 12053
rect 36078 12044 36084 12056
rect 36136 12044 36142 12096
rect 36173 12087 36231 12093
rect 36173 12053 36185 12087
rect 36219 12084 36231 12087
rect 36814 12084 36820 12096
rect 36219 12056 36820 12084
rect 36219 12053 36231 12056
rect 36173 12047 36231 12053
rect 36814 12044 36820 12056
rect 36872 12044 36878 12096
rect 1104 11994 39352 12016
rect 1104 11942 10472 11994
rect 10524 11942 10536 11994
rect 10588 11942 10600 11994
rect 10652 11942 10664 11994
rect 10716 11942 10728 11994
rect 10780 11942 19994 11994
rect 20046 11942 20058 11994
rect 20110 11942 20122 11994
rect 20174 11942 20186 11994
rect 20238 11942 20250 11994
rect 20302 11942 29516 11994
rect 29568 11942 29580 11994
rect 29632 11942 29644 11994
rect 29696 11942 29708 11994
rect 29760 11942 29772 11994
rect 29824 11942 39038 11994
rect 39090 11942 39102 11994
rect 39154 11942 39166 11994
rect 39218 11942 39230 11994
rect 39282 11942 39294 11994
rect 39346 11942 39352 11994
rect 1104 11920 39352 11942
rect 2222 11840 2228 11892
rect 2280 11880 2286 11892
rect 2866 11880 2872 11892
rect 2280 11852 2872 11880
rect 2280 11840 2286 11852
rect 1762 11704 1768 11756
rect 1820 11704 1826 11756
rect 2424 11753 2452 11852
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 3418 11840 3424 11892
rect 3476 11880 3482 11892
rect 5350 11880 5356 11892
rect 3476 11852 5356 11880
rect 3476 11840 3482 11852
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 5500 11852 6561 11880
rect 5500 11840 5506 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 6549 11843 6607 11849
rect 6638 11840 6644 11892
rect 6696 11880 6702 11892
rect 7193 11883 7251 11889
rect 7193 11880 7205 11883
rect 6696 11852 7205 11880
rect 6696 11840 6702 11852
rect 7193 11849 7205 11852
rect 7239 11849 7251 11883
rect 7193 11843 7251 11849
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 7892 11852 9168 11880
rect 7892 11840 7898 11852
rect 6454 11812 6460 11824
rect 4816 11784 6460 11812
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11713 2467 11747
rect 2409 11707 2467 11713
rect 3786 11704 3792 11756
rect 3844 11704 3850 11756
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 4816 11676 4844 11784
rect 6454 11772 6460 11784
rect 6512 11772 6518 11824
rect 6822 11772 6828 11824
rect 6880 11812 6886 11824
rect 9140 11812 9168 11852
rect 9306 11840 9312 11892
rect 9364 11880 9370 11892
rect 9766 11880 9772 11892
rect 9364 11852 9772 11880
rect 9364 11840 9370 11852
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10962 11880 10968 11892
rect 10244 11852 10968 11880
rect 10244 11812 10272 11852
rect 6880 11784 9076 11812
rect 9140 11784 10272 11812
rect 6880 11772 6886 11784
rect 5626 11704 5632 11756
rect 5684 11704 5690 11756
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 7006 11744 7012 11756
rect 6963 11716 7012 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 2731 11648 4844 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 5736 11676 5764 11707
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 7282 11704 7288 11756
rect 7340 11704 7346 11756
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 7984 11716 8033 11744
rect 7984 11704 7990 11716
rect 8021 11713 8033 11716
rect 8067 11713 8079 11747
rect 8205 11747 8263 11753
rect 8205 11744 8217 11747
rect 8021 11707 8079 11713
rect 8128 11716 8217 11744
rect 8128 11688 8156 11716
rect 8205 11713 8217 11716
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 9048 11753 9076 11784
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11713 8447 11747
rect 8389 11707 8447 11713
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11744 9091 11747
rect 9858 11744 9864 11756
rect 9079 11716 9864 11744
rect 9079 11713 9091 11716
rect 9033 11707 9091 11713
rect 5592 11648 5764 11676
rect 5592 11636 5598 11648
rect 5810 11636 5816 11688
rect 5868 11636 5874 11688
rect 7374 11676 7380 11688
rect 6840 11648 7380 11676
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 6840 11608 6868 11648
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 8110 11636 8116 11688
rect 8168 11636 8174 11688
rect 8404 11676 8432 11707
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11744 10103 11747
rect 10778 11744 10784 11756
rect 10091 11716 10784 11744
rect 10091 11713 10103 11716
rect 10045 11707 10103 11713
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 10137 11679 10195 11685
rect 8220 11648 9996 11676
rect 4203 11580 6868 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 7742 11568 7748 11620
rect 7800 11608 7806 11620
rect 8220 11608 8248 11648
rect 7800 11580 8248 11608
rect 7800 11568 7806 11580
rect 8478 11568 8484 11620
rect 8536 11608 8542 11620
rect 8573 11611 8631 11617
rect 8573 11608 8585 11611
rect 8536 11580 8585 11608
rect 8536 11568 8542 11580
rect 8573 11577 8585 11580
rect 8619 11577 8631 11611
rect 8573 11571 8631 11577
rect 9125 11611 9183 11617
rect 9125 11577 9137 11611
rect 9171 11608 9183 11611
rect 9582 11608 9588 11620
rect 9171 11580 9588 11608
rect 9171 11577 9183 11580
rect 9125 11571 9183 11577
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 1854 11500 1860 11552
rect 1912 11500 1918 11552
rect 2038 11500 2044 11552
rect 2096 11540 2102 11552
rect 2682 11540 2688 11552
rect 2096 11512 2688 11540
rect 2096 11500 2102 11512
rect 2682 11500 2688 11512
rect 2740 11500 2746 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 5261 11543 5319 11549
rect 5261 11540 5273 11543
rect 4304 11512 5273 11540
rect 4304 11500 4310 11512
rect 5261 11509 5273 11512
rect 5307 11509 5319 11543
rect 5261 11503 5319 11509
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6328 11512 6837 11540
rect 6328 11500 6334 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 7006 11500 7012 11552
rect 7064 11500 7070 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 9456 11512 9689 11540
rect 9456 11500 9462 11512
rect 9677 11509 9689 11512
rect 9723 11509 9735 11543
rect 9968 11540 9996 11648
rect 10137 11645 10149 11679
rect 10183 11645 10195 11679
rect 10137 11639 10195 11645
rect 10152 11608 10180 11639
rect 10318 11636 10324 11688
rect 10376 11636 10382 11688
rect 10888 11676 10916 11852
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 13814 11880 13820 11892
rect 12406 11852 13820 11880
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11744 11023 11747
rect 11238 11744 11244 11756
rect 11011 11716 11244 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 11238 11704 11244 11716
rect 11296 11744 11302 11756
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 11296 11716 12265 11744
rect 11296 11704 11302 11716
rect 12253 11713 12265 11716
rect 12299 11744 12311 11747
rect 12406 11744 12434 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 13906 11840 13912 11892
rect 13964 11880 13970 11892
rect 15654 11880 15660 11892
rect 13964 11852 15660 11880
rect 13964 11840 13970 11852
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 16301 11883 16359 11889
rect 16301 11849 16313 11883
rect 16347 11880 16359 11883
rect 16850 11880 16856 11892
rect 16347 11852 16856 11880
rect 16347 11849 16359 11852
rect 16301 11843 16359 11849
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 17954 11880 17960 11892
rect 16960 11852 17960 11880
rect 13170 11772 13176 11824
rect 13228 11772 13234 11824
rect 15838 11812 15844 11824
rect 14398 11784 15844 11812
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 12299 11716 12434 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12676 11716 12909 11744
rect 12676 11704 12682 11716
rect 12897 11713 12909 11716
rect 12943 11713 12955 11747
rect 16022 11744 16028 11756
rect 12897 11707 12955 11713
rect 14844 11716 16028 11744
rect 14844 11676 14872 11716
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16960 11744 16988 11852
rect 17954 11840 17960 11852
rect 18012 11880 18018 11892
rect 18690 11880 18696 11892
rect 18012 11852 18696 11880
rect 18012 11840 18018 11852
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 18966 11840 18972 11892
rect 19024 11880 19030 11892
rect 19521 11883 19579 11889
rect 19521 11880 19533 11883
rect 19024 11852 19533 11880
rect 19024 11840 19030 11852
rect 19521 11849 19533 11852
rect 19567 11849 19579 11883
rect 19521 11843 19579 11849
rect 20073 11883 20131 11889
rect 20073 11849 20085 11883
rect 20119 11849 20131 11883
rect 20073 11843 20131 11849
rect 17494 11772 17500 11824
rect 17552 11772 17558 11824
rect 18506 11772 18512 11824
rect 18564 11812 18570 11824
rect 20088 11812 20116 11843
rect 20438 11840 20444 11892
rect 20496 11840 20502 11892
rect 20530 11840 20536 11892
rect 20588 11840 20594 11892
rect 22370 11880 22376 11892
rect 21100 11852 22376 11880
rect 21100 11812 21128 11852
rect 22370 11840 22376 11852
rect 22428 11840 22434 11892
rect 25130 11880 25136 11892
rect 23216 11852 25136 11880
rect 21818 11812 21824 11824
rect 18564 11784 18828 11812
rect 20088 11784 21128 11812
rect 21192 11784 21824 11812
rect 18564 11772 18570 11784
rect 16163 11716 16988 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 17092 11716 17141 11744
rect 17092 11704 17098 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17277 11747 17335 11753
rect 17277 11713 17289 11747
rect 17323 11713 17335 11747
rect 17277 11707 17335 11713
rect 10888 11648 14872 11676
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11676 15991 11679
rect 16206 11676 16212 11688
rect 15979 11648 16212 11676
rect 15979 11645 15991 11648
rect 15933 11639 15991 11645
rect 10410 11608 10416 11620
rect 10152 11580 10416 11608
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 12434 11608 12440 11620
rect 10520 11580 12440 11608
rect 10520 11540 10548 11580
rect 12434 11568 12440 11580
rect 12492 11568 12498 11620
rect 14936 11608 14964 11639
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 16298 11636 16304 11688
rect 16356 11676 16362 11688
rect 17292 11676 17320 11707
rect 17402 11704 17408 11756
rect 17460 11704 17466 11756
rect 17635 11747 17693 11753
rect 17635 11713 17647 11747
rect 17681 11744 17693 11747
rect 17862 11744 17868 11756
rect 17681 11716 17868 11744
rect 17681 11713 17693 11716
rect 17635 11707 17693 11713
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18230 11744 18236 11756
rect 18012 11716 18236 11744
rect 18012 11704 18018 11716
rect 18230 11704 18236 11716
rect 18288 11704 18294 11756
rect 18598 11704 18604 11756
rect 18656 11704 18662 11756
rect 18800 11685 18828 11784
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11744 19487 11747
rect 19518 11744 19524 11756
rect 19475 11716 19524 11744
rect 19475 11713 19487 11716
rect 19429 11707 19487 11713
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 21192 11744 21220 11784
rect 21818 11772 21824 11784
rect 21876 11772 21882 11824
rect 22094 11772 22100 11824
rect 22152 11812 22158 11824
rect 22281 11815 22339 11821
rect 22281 11812 22293 11815
rect 22152 11784 22293 11812
rect 22152 11772 22158 11784
rect 22281 11781 22293 11784
rect 22327 11781 22339 11815
rect 22281 11775 22339 11781
rect 22922 11772 22928 11824
rect 22980 11812 22986 11824
rect 23216 11812 23244 11852
rect 25130 11840 25136 11852
rect 25188 11840 25194 11892
rect 25317 11883 25375 11889
rect 25317 11849 25329 11883
rect 25363 11849 25375 11883
rect 25317 11843 25375 11849
rect 22980 11784 23244 11812
rect 22980 11772 22986 11784
rect 20496 11716 21220 11744
rect 21269 11747 21327 11753
rect 20496 11704 20502 11716
rect 21269 11713 21281 11747
rect 21315 11744 21327 11747
rect 21634 11744 21640 11756
rect 21315 11716 21640 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 21634 11704 21640 11716
rect 21692 11704 21698 11756
rect 21726 11704 21732 11756
rect 21784 11744 21790 11756
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 21784 11716 22017 11744
rect 21784 11704 21790 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 22373 11747 22431 11753
rect 22373 11713 22385 11747
rect 22419 11744 22431 11747
rect 22646 11744 22652 11756
rect 22419 11716 22652 11744
rect 22419 11713 22431 11716
rect 22373 11707 22431 11713
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 16356 11648 18705 11676
rect 16356 11636 16362 11648
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 18785 11679 18843 11685
rect 18785 11645 18797 11679
rect 18831 11645 18843 11679
rect 18785 11639 18843 11645
rect 19702 11636 19708 11688
rect 19760 11676 19766 11688
rect 20625 11679 20683 11685
rect 20625 11676 20637 11679
rect 19760 11648 20637 11676
rect 19760 11636 19766 11648
rect 20625 11645 20637 11648
rect 20671 11645 20683 11679
rect 22204 11676 22232 11707
rect 22646 11704 22652 11716
rect 22704 11704 22710 11756
rect 23124 11753 23152 11784
rect 23934 11772 23940 11824
rect 23992 11772 23998 11824
rect 24762 11772 24768 11824
rect 24820 11812 24826 11824
rect 25332 11812 25360 11843
rect 26050 11840 26056 11892
rect 26108 11880 26114 11892
rect 26108 11852 28764 11880
rect 26108 11840 26114 11852
rect 24820 11784 25360 11812
rect 25685 11815 25743 11821
rect 24820 11772 24826 11784
rect 25685 11781 25697 11815
rect 25731 11812 25743 11815
rect 25774 11812 25780 11824
rect 25731 11784 25780 11812
rect 25731 11781 25743 11784
rect 25685 11775 25743 11781
rect 25774 11772 25780 11784
rect 25832 11772 25838 11824
rect 26418 11812 26424 11824
rect 25884 11784 26424 11812
rect 23109 11747 23167 11753
rect 23109 11713 23121 11747
rect 23155 11713 23167 11747
rect 25884 11744 25912 11784
rect 26418 11772 26424 11784
rect 26476 11772 26482 11824
rect 27433 11815 27491 11821
rect 27433 11781 27445 11815
rect 27479 11812 27491 11815
rect 27522 11812 27528 11824
rect 27479 11784 27528 11812
rect 27479 11781 27491 11784
rect 27433 11775 27491 11781
rect 27522 11772 27528 11784
rect 27580 11772 27586 11824
rect 28166 11772 28172 11824
rect 28224 11772 28230 11824
rect 23109 11707 23167 11713
rect 25792 11716 25912 11744
rect 22204 11648 22416 11676
rect 20625 11639 20683 11645
rect 22388 11620 22416 11648
rect 22462 11636 22468 11688
rect 22520 11676 22526 11688
rect 25792 11685 25820 11716
rect 25958 11704 25964 11756
rect 26016 11744 26022 11756
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 26016 11716 27169 11744
rect 26016 11704 26022 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 28736 11744 28764 11852
rect 28902 11840 28908 11892
rect 28960 11840 28966 11892
rect 29178 11840 29184 11892
rect 29236 11880 29242 11892
rect 31113 11883 31171 11889
rect 31113 11880 31125 11883
rect 29236 11852 31125 11880
rect 29236 11840 29242 11852
rect 31113 11849 31125 11852
rect 31159 11849 31171 11883
rect 31113 11843 31171 11849
rect 32677 11883 32735 11889
rect 32677 11849 32689 11883
rect 32723 11849 32735 11883
rect 32677 11843 32735 11849
rect 33045 11883 33103 11889
rect 33045 11849 33057 11883
rect 33091 11880 33103 11883
rect 33410 11880 33416 11892
rect 33091 11852 33416 11880
rect 33091 11849 33103 11852
rect 33045 11843 33103 11849
rect 29454 11772 29460 11824
rect 29512 11772 29518 11824
rect 29657 11815 29715 11821
rect 29657 11812 29669 11815
rect 29564 11784 29669 11812
rect 29564 11744 29592 11784
rect 29657 11781 29669 11784
rect 29703 11781 29715 11815
rect 29657 11775 29715 11781
rect 30006 11772 30012 11824
rect 30064 11812 30070 11824
rect 31754 11812 31760 11824
rect 30064 11784 31760 11812
rect 30064 11772 30070 11784
rect 31754 11772 31760 11784
rect 31812 11812 31818 11824
rect 32306 11812 32312 11824
rect 31812 11784 32312 11812
rect 31812 11772 31818 11784
rect 32306 11772 32312 11784
rect 32364 11772 32370 11824
rect 32692 11812 32720 11843
rect 33410 11840 33416 11852
rect 33468 11880 33474 11892
rect 36633 11883 36691 11889
rect 36633 11880 36645 11883
rect 33468 11852 36645 11880
rect 33468 11840 33474 11852
rect 36633 11849 36645 11852
rect 36679 11849 36691 11883
rect 36633 11843 36691 11849
rect 35161 11815 35219 11821
rect 35161 11812 35173 11815
rect 32692 11784 35173 11812
rect 35161 11781 35173 11784
rect 35207 11781 35219 11815
rect 38105 11815 38163 11821
rect 38105 11812 38117 11815
rect 36386 11784 38117 11812
rect 35161 11775 35219 11781
rect 38105 11781 38117 11784
rect 38151 11781 38163 11815
rect 38105 11775 38163 11781
rect 30558 11744 30564 11756
rect 28736 11716 30564 11744
rect 27157 11707 27215 11713
rect 30558 11704 30564 11716
rect 30616 11704 30622 11756
rect 30742 11704 30748 11756
rect 30800 11744 30806 11756
rect 30929 11747 30987 11753
rect 30929 11744 30941 11747
rect 30800 11716 30941 11744
rect 30800 11704 30806 11716
rect 30929 11713 30941 11716
rect 30975 11713 30987 11747
rect 30929 11707 30987 11713
rect 31386 11704 31392 11756
rect 31444 11744 31450 11756
rect 31444 11716 32352 11744
rect 31444 11704 31450 11716
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 22520 11648 23397 11676
rect 22520 11636 22526 11648
rect 23385 11645 23397 11648
rect 23431 11645 23443 11679
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 23385 11639 23443 11645
rect 24412 11648 25789 11676
rect 14936 11580 22324 11608
rect 9968 11512 10548 11540
rect 9677 11503 9735 11509
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 10928 11512 11069 11540
rect 10928 11500 10934 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 11057 11503 11115 11509
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 12345 11543 12403 11549
rect 12345 11540 12357 11543
rect 12308 11512 12357 11540
rect 12308 11500 12314 11512
rect 12345 11509 12357 11512
rect 12391 11509 12403 11543
rect 12345 11503 12403 11509
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13722 11540 13728 11552
rect 13044 11512 13728 11540
rect 13044 11500 13050 11512
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 14458 11500 14464 11552
rect 14516 11540 14522 11552
rect 15654 11540 15660 11552
rect 14516 11512 15660 11540
rect 14516 11500 14522 11512
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 16724 11512 17785 11540
rect 16724 11500 16730 11512
rect 17773 11509 17785 11512
rect 17819 11509 17831 11543
rect 17773 11503 17831 11509
rect 18230 11500 18236 11552
rect 18288 11500 18294 11552
rect 18414 11500 18420 11552
rect 18472 11540 18478 11552
rect 20714 11540 20720 11552
rect 18472 11512 20720 11540
rect 18472 11500 18478 11512
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 21358 11500 21364 11552
rect 21416 11500 21422 11552
rect 22296 11540 22324 11580
rect 22370 11568 22376 11620
rect 22428 11568 22434 11620
rect 22480 11580 23244 11608
rect 22480 11540 22508 11580
rect 22296 11512 22508 11540
rect 22554 11500 22560 11552
rect 22612 11500 22618 11552
rect 23216 11540 23244 11580
rect 24412 11540 24440 11648
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 25869 11679 25927 11685
rect 25869 11645 25881 11679
rect 25915 11676 25927 11679
rect 26142 11676 26148 11688
rect 25915 11648 26148 11676
rect 25915 11645 25927 11648
rect 25869 11639 25927 11645
rect 25590 11568 25596 11620
rect 25648 11608 25654 11620
rect 25884 11608 25912 11639
rect 26142 11636 26148 11648
rect 26200 11636 26206 11688
rect 27890 11636 27896 11688
rect 27948 11676 27954 11688
rect 29086 11676 29092 11688
rect 27948 11648 29092 11676
rect 27948 11636 27954 11648
rect 29086 11636 29092 11648
rect 29144 11636 29150 11688
rect 30469 11679 30527 11685
rect 30469 11645 30481 11679
rect 30515 11676 30527 11679
rect 31110 11676 31116 11688
rect 30515 11648 31116 11676
rect 30515 11645 30527 11648
rect 30469 11639 30527 11645
rect 31110 11636 31116 11648
rect 31168 11636 31174 11688
rect 31202 11636 31208 11688
rect 31260 11676 31266 11688
rect 32122 11676 32128 11688
rect 31260 11648 32128 11676
rect 31260 11636 31266 11648
rect 32122 11636 32128 11648
rect 32180 11636 32186 11688
rect 32324 11676 32352 11716
rect 32398 11704 32404 11756
rect 32456 11744 32462 11756
rect 33042 11744 33048 11756
rect 32456 11716 33048 11744
rect 32456 11704 32462 11716
rect 33042 11704 33048 11716
rect 33100 11744 33106 11756
rect 33873 11747 33931 11753
rect 33100 11716 33272 11744
rect 33100 11704 33106 11716
rect 32582 11676 32588 11688
rect 32324 11648 32588 11676
rect 32582 11636 32588 11648
rect 32640 11636 32646 11688
rect 33134 11636 33140 11688
rect 33192 11636 33198 11688
rect 33244 11685 33272 11716
rect 33873 11713 33885 11747
rect 33919 11744 33931 11747
rect 33962 11744 33968 11756
rect 33919 11716 33968 11744
rect 33919 11713 33931 11716
rect 33873 11707 33931 11713
rect 33962 11704 33968 11716
rect 34020 11744 34026 11756
rect 34790 11744 34796 11756
rect 34020 11716 34796 11744
rect 34020 11704 34026 11716
rect 34790 11704 34796 11716
rect 34848 11704 34854 11756
rect 38010 11704 38016 11756
rect 38068 11704 38074 11756
rect 33229 11679 33287 11685
rect 33229 11645 33241 11679
rect 33275 11645 33287 11679
rect 33229 11639 33287 11645
rect 34606 11636 34612 11688
rect 34664 11676 34670 11688
rect 34885 11679 34943 11685
rect 34885 11676 34897 11679
rect 34664 11648 34897 11676
rect 34664 11636 34670 11648
rect 34885 11645 34897 11648
rect 34931 11645 34943 11679
rect 35894 11676 35900 11688
rect 34885 11639 34943 11645
rect 34992 11648 35900 11676
rect 25648 11580 25912 11608
rect 25648 11568 25654 11580
rect 26234 11568 26240 11620
rect 26292 11608 26298 11620
rect 26878 11608 26884 11620
rect 26292 11580 26884 11608
rect 26292 11568 26298 11580
rect 26878 11568 26884 11580
rect 26936 11568 26942 11620
rect 28718 11568 28724 11620
rect 28776 11608 28782 11620
rect 29825 11611 29883 11617
rect 28776 11580 29684 11608
rect 28776 11568 28782 11580
rect 29656 11552 29684 11580
rect 29825 11577 29837 11611
rect 29871 11608 29883 11611
rect 30745 11611 30803 11617
rect 30745 11608 30757 11611
rect 29871 11580 30757 11608
rect 29871 11577 29883 11580
rect 29825 11571 29883 11577
rect 30745 11577 30757 11580
rect 30791 11577 30803 11611
rect 30745 11571 30803 11577
rect 30837 11611 30895 11617
rect 30837 11577 30849 11611
rect 30883 11608 30895 11611
rect 33318 11608 33324 11620
rect 30883 11580 33324 11608
rect 30883 11577 30895 11580
rect 30837 11571 30895 11577
rect 33318 11568 33324 11580
rect 33376 11568 33382 11620
rect 34992 11608 35020 11648
rect 35894 11636 35900 11648
rect 35952 11636 35958 11688
rect 33796 11580 35020 11608
rect 23216 11512 24440 11540
rect 24857 11543 24915 11549
rect 24857 11509 24869 11543
rect 24903 11540 24915 11543
rect 25130 11540 25136 11552
rect 24903 11512 25136 11540
rect 24903 11509 24915 11512
rect 24857 11503 24915 11509
rect 25130 11500 25136 11512
rect 25188 11500 25194 11552
rect 25682 11500 25688 11552
rect 25740 11540 25746 11552
rect 29362 11540 29368 11552
rect 25740 11512 29368 11540
rect 25740 11500 25746 11512
rect 29362 11500 29368 11512
rect 29420 11500 29426 11552
rect 29638 11500 29644 11552
rect 29696 11500 29702 11552
rect 30558 11500 30564 11552
rect 30616 11540 30622 11552
rect 33796 11540 33824 11580
rect 30616 11512 33824 11540
rect 30616 11500 30622 11512
rect 33962 11500 33968 11552
rect 34020 11500 34026 11552
rect 1104 11450 39192 11472
rect 1104 11398 5711 11450
rect 5763 11398 5775 11450
rect 5827 11398 5839 11450
rect 5891 11398 5903 11450
rect 5955 11398 5967 11450
rect 6019 11398 15233 11450
rect 15285 11398 15297 11450
rect 15349 11398 15361 11450
rect 15413 11398 15425 11450
rect 15477 11398 15489 11450
rect 15541 11398 24755 11450
rect 24807 11398 24819 11450
rect 24871 11398 24883 11450
rect 24935 11398 24947 11450
rect 24999 11398 25011 11450
rect 25063 11398 34277 11450
rect 34329 11398 34341 11450
rect 34393 11398 34405 11450
rect 34457 11398 34469 11450
rect 34521 11398 34533 11450
rect 34585 11398 39192 11450
rect 1104 11376 39192 11398
rect 2685 11339 2743 11345
rect 2685 11305 2697 11339
rect 2731 11336 2743 11339
rect 3878 11336 3884 11348
rect 2731 11308 3884 11336
rect 2731 11305 2743 11308
rect 2685 11299 2743 11305
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 4396 11308 7941 11336
rect 4396 11296 4402 11308
rect 7929 11305 7941 11308
rect 7975 11305 7987 11339
rect 7929 11299 7987 11305
rect 8478 11296 8484 11348
rect 8536 11296 8542 11348
rect 9122 11336 9128 11348
rect 8588 11308 9128 11336
rect 3050 11228 3056 11280
rect 3108 11268 3114 11280
rect 3108 11240 4108 11268
rect 3108 11228 3114 11240
rect 3142 11160 3148 11212
rect 3200 11160 3206 11212
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11200 3387 11203
rect 3418 11200 3424 11212
rect 3375 11172 3424 11200
rect 3375 11169 3387 11172
rect 3329 11163 3387 11169
rect 3418 11160 3424 11172
rect 3476 11160 3482 11212
rect 4080 11200 4108 11240
rect 5350 11228 5356 11280
rect 5408 11268 5414 11280
rect 5408 11240 5948 11268
rect 5408 11228 5414 11240
rect 5626 11200 5632 11212
rect 4080 11172 5632 11200
rect 5626 11160 5632 11172
rect 5684 11200 5690 11212
rect 5721 11203 5779 11209
rect 5721 11200 5733 11203
rect 5684 11172 5733 11200
rect 5684 11160 5690 11172
rect 5721 11169 5733 11172
rect 5767 11169 5779 11203
rect 5721 11163 5779 11169
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2087 11104 2774 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 934 11024 940 11076
rect 992 11064 998 11076
rect 1673 11067 1731 11073
rect 1673 11064 1685 11067
rect 992 11036 1685 11064
rect 992 11024 998 11036
rect 1673 11033 1685 11036
rect 1719 11033 1731 11067
rect 1673 11027 1731 11033
rect 2746 10996 2774 11104
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 3970 11132 3976 11144
rect 2924 11104 3976 11132
rect 2924 11092 2930 11104
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 5920 11132 5948 11240
rect 5994 11228 6000 11280
rect 6052 11268 6058 11280
rect 6270 11268 6276 11280
rect 6052 11240 6276 11268
rect 6052 11228 6058 11240
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 6365 11271 6423 11277
rect 6365 11237 6377 11271
rect 6411 11268 6423 11271
rect 8110 11268 8116 11280
rect 6411 11240 8116 11268
rect 6411 11237 6423 11240
rect 6365 11231 6423 11237
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 8294 11228 8300 11280
rect 8352 11268 8358 11280
rect 8588 11268 8616 11308
rect 9122 11296 9128 11308
rect 9180 11336 9186 11348
rect 9180 11308 10456 11336
rect 9180 11296 9186 11308
rect 8352 11240 8616 11268
rect 10428 11268 10456 11308
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10560 11308 10885 11336
rect 10560 11296 10566 11308
rect 10873 11305 10885 11308
rect 10919 11336 10931 11339
rect 11606 11336 11612 11348
rect 10919 11308 11612 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 15654 11336 15660 11348
rect 12492 11308 15660 11336
rect 12492 11296 12498 11308
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16117 11339 16175 11345
rect 16117 11305 16129 11339
rect 16163 11336 16175 11339
rect 16298 11336 16304 11348
rect 16163 11308 16304 11336
rect 16163 11305 16175 11308
rect 16117 11299 16175 11305
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 17126 11296 17132 11348
rect 17184 11336 17190 11348
rect 17310 11336 17316 11348
rect 17184 11308 17316 11336
rect 17184 11296 17190 11308
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 17494 11296 17500 11348
rect 17552 11336 17558 11348
rect 17552 11308 18368 11336
rect 17552 11296 17558 11308
rect 13630 11268 13636 11280
rect 10428 11240 13636 11268
rect 8352 11228 8358 11240
rect 13630 11228 13636 11240
rect 13688 11228 13694 11280
rect 18230 11268 18236 11280
rect 15764 11240 18236 11268
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 7708 11172 9137 11200
rect 7708 11160 7714 11172
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 9398 11160 9404 11212
rect 9456 11160 9462 11212
rect 11882 11160 11888 11212
rect 11940 11160 11946 11212
rect 12618 11160 12624 11212
rect 12676 11200 12682 11212
rect 14369 11203 14427 11209
rect 14369 11200 14381 11203
rect 12676 11172 14381 11200
rect 12676 11160 12682 11172
rect 14369 11169 14381 11172
rect 14415 11169 14427 11203
rect 14369 11163 14427 11169
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11200 14703 11203
rect 15764 11200 15792 11240
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 18340 11268 18368 11308
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 19610 11336 19616 11348
rect 18472 11308 19616 11336
rect 18472 11296 18478 11308
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 21634 11336 21640 11348
rect 20088 11308 21640 11336
rect 18340 11240 18644 11268
rect 14691 11172 15792 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 16022 11160 16028 11212
rect 16080 11200 16086 11212
rect 17313 11203 17371 11209
rect 17313 11200 17325 11203
rect 16080 11172 17325 11200
rect 16080 11160 16086 11172
rect 17313 11169 17325 11172
rect 17359 11200 17371 11203
rect 17402 11200 17408 11212
rect 17359 11172 17408 11200
rect 17359 11169 17371 11172
rect 17313 11163 17371 11169
rect 17402 11160 17408 11172
rect 17460 11200 17466 11212
rect 18509 11203 18567 11209
rect 18509 11200 18521 11203
rect 17460 11172 18521 11200
rect 17460 11160 17466 11172
rect 18509 11169 18521 11172
rect 18555 11169 18567 11203
rect 18616 11200 18644 11240
rect 18616 11172 19334 11200
rect 18509 11163 18567 11169
rect 6270 11132 6276 11144
rect 5920 11104 6276 11132
rect 6270 11092 6276 11104
rect 6328 11132 6334 11144
rect 6822 11132 6828 11144
rect 6328 11104 6828 11132
rect 6328 11092 6334 11104
rect 6822 11092 6828 11104
rect 6880 11132 6886 11144
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6880 11104 6929 11132
rect 6880 11092 6886 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7524 11104 7573 11132
rect 7524 11092 7530 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 7742 11092 7748 11144
rect 7800 11092 7806 11144
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11132 8447 11135
rect 8478 11132 8484 11144
rect 8435 11104 8484 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 8478 11092 8484 11104
rect 8536 11132 8542 11144
rect 8938 11132 8944 11144
rect 8536 11104 8944 11132
rect 8536 11092 8542 11104
rect 8938 11092 8944 11104
rect 8996 11092 9002 11144
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11132 11759 11135
rect 11790 11132 11796 11144
rect 11747 11104 11796 11132
rect 11747 11101 11759 11104
rect 11701 11095 11759 11101
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 13538 11132 13544 11144
rect 12032 11104 13544 11132
rect 12032 11092 12038 11104
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 18012 11104 18245 11132
rect 18012 11092 18018 11104
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 19306 11132 19334 11172
rect 19429 11135 19487 11141
rect 19429 11132 19441 11135
rect 19306 11104 19441 11132
rect 18233 11095 18291 11101
rect 19429 11101 19441 11104
rect 19475 11132 19487 11135
rect 20088 11132 20116 11308
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 21729 11339 21787 11345
rect 21729 11305 21741 11339
rect 21775 11336 21787 11339
rect 21818 11336 21824 11348
rect 21775 11308 21824 11336
rect 21775 11305 21787 11308
rect 21729 11299 21787 11305
rect 21818 11296 21824 11308
rect 21876 11296 21882 11348
rect 22646 11336 22652 11348
rect 22066 11308 22652 11336
rect 20165 11271 20223 11277
rect 20165 11237 20177 11271
rect 20211 11268 20223 11271
rect 22066 11268 22094 11308
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 23934 11296 23940 11348
rect 23992 11296 23998 11348
rect 25590 11336 25596 11348
rect 25240 11308 25596 11336
rect 25130 11268 25136 11280
rect 20211 11240 22094 11268
rect 22204 11240 25136 11268
rect 20211 11237 20223 11240
rect 20165 11231 20223 11237
rect 20714 11160 20720 11212
rect 20772 11160 20778 11212
rect 22204 11209 22232 11240
rect 25130 11228 25136 11240
rect 25188 11228 25194 11280
rect 22189 11203 22247 11209
rect 22189 11169 22201 11203
rect 22235 11169 22247 11203
rect 22189 11163 22247 11169
rect 22373 11203 22431 11209
rect 22373 11169 22385 11203
rect 22419 11200 22431 11203
rect 25240 11200 25268 11308
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 26326 11296 26332 11348
rect 26384 11336 26390 11348
rect 26384 11308 26556 11336
rect 26384 11296 26390 11308
rect 25682 11268 25688 11280
rect 22419 11172 25268 11200
rect 25332 11240 25688 11268
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 19475 11104 20116 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 20530 11092 20536 11144
rect 20588 11132 20594 11144
rect 23750 11132 23756 11144
rect 20588 11104 23756 11132
rect 20588 11092 20594 11104
rect 23750 11092 23756 11104
rect 23808 11092 23814 11144
rect 23842 11092 23848 11144
rect 23900 11132 23906 11144
rect 24578 11132 24584 11144
rect 23900 11104 24584 11132
rect 23900 11092 23906 11104
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 25332 11132 25360 11240
rect 25682 11228 25688 11240
rect 25740 11228 25746 11280
rect 25777 11203 25835 11209
rect 25777 11169 25789 11203
rect 25823 11200 25835 11203
rect 26050 11200 26056 11212
rect 25823 11172 26056 11200
rect 25823 11169 25835 11172
rect 25777 11163 25835 11169
rect 26050 11160 26056 11172
rect 26108 11160 26114 11212
rect 26418 11160 26424 11212
rect 26476 11160 26482 11212
rect 24688 11104 25360 11132
rect 25501 11135 25559 11141
rect 3053 11067 3111 11073
rect 3053 11033 3065 11067
rect 3099 11064 3111 11067
rect 3878 11064 3884 11076
rect 3099 11036 3884 11064
rect 3099 11033 3111 11036
rect 3053 11027 3111 11033
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4246 11024 4252 11076
rect 4304 11024 4310 11076
rect 5626 11064 5632 11076
rect 5474 11036 5632 11064
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 7009 11067 7067 11073
rect 7009 11033 7021 11067
rect 7055 11064 7067 11067
rect 13633 11067 13691 11073
rect 7055 11036 9890 11064
rect 7055 11033 7067 11036
rect 7009 11027 7067 11033
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 13679 11036 14596 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 6086 10996 6092 11008
rect 2746 10968 6092 10996
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 9306 10996 9312 11008
rect 6880 10968 9312 10996
rect 6880 10956 6886 10968
rect 9306 10956 9312 10968
rect 9364 10956 9370 11008
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 11882 10996 11888 11008
rect 10284 10968 11888 10996
rect 10284 10956 10290 10968
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 14568 10996 14596 11036
rect 14752 11036 15134 11064
rect 14752 10996 14780 11036
rect 16206 11024 16212 11076
rect 16264 11064 16270 11076
rect 17221 11067 17279 11073
rect 17221 11064 17233 11067
rect 16264 11036 17233 11064
rect 16264 11024 16270 11036
rect 17221 11033 17233 11036
rect 17267 11064 17279 11067
rect 18506 11064 18512 11076
rect 17267 11036 18512 11064
rect 17267 11033 17279 11036
rect 17221 11027 17279 11033
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 20625 11067 20683 11073
rect 20625 11064 20637 11067
rect 19444 11036 20637 11064
rect 19444 11008 19472 11036
rect 20625 11033 20637 11036
rect 20671 11033 20683 11067
rect 20625 11027 20683 11033
rect 23014 11024 23020 11076
rect 23072 11024 23078 11076
rect 23201 11067 23259 11073
rect 23201 11033 23213 11067
rect 23247 11064 23259 11067
rect 23566 11064 23572 11076
rect 23247 11036 23572 11064
rect 23247 11033 23259 11036
rect 23201 11027 23259 11033
rect 23566 11024 23572 11036
rect 23624 11024 23630 11076
rect 24302 11024 24308 11076
rect 24360 11064 24366 11076
rect 24688 11064 24716 11104
rect 25501 11101 25513 11135
rect 25547 11132 25559 11135
rect 26234 11132 26240 11144
rect 25547 11104 26240 11132
rect 25547 11101 25559 11104
rect 25501 11095 25559 11101
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 26329 11135 26387 11141
rect 26329 11101 26341 11135
rect 26375 11132 26387 11135
rect 26436 11132 26464 11160
rect 26528 11141 26556 11308
rect 26602 11296 26608 11348
rect 26660 11296 26666 11348
rect 28258 11296 28264 11348
rect 28316 11336 28322 11348
rect 29270 11336 29276 11348
rect 28316 11308 29276 11336
rect 28316 11296 28322 11308
rect 29270 11296 29276 11308
rect 29328 11336 29334 11348
rect 29454 11336 29460 11348
rect 29328 11308 29460 11336
rect 29328 11296 29334 11308
rect 29454 11296 29460 11308
rect 29512 11296 29518 11348
rect 30745 11339 30803 11345
rect 30745 11305 30757 11339
rect 30791 11336 30803 11339
rect 31294 11336 31300 11348
rect 30791 11308 31300 11336
rect 30791 11305 30803 11308
rect 30745 11299 30803 11305
rect 31294 11296 31300 11308
rect 31352 11296 31358 11348
rect 34974 11296 34980 11348
rect 35032 11296 35038 11348
rect 36078 11296 36084 11348
rect 36136 11336 36142 11348
rect 36265 11339 36323 11345
rect 36265 11336 36277 11339
rect 36136 11308 36277 11336
rect 36136 11296 36142 11308
rect 36265 11305 36277 11308
rect 36311 11305 36323 11339
rect 36265 11299 36323 11305
rect 26620 11268 26648 11296
rect 27154 11268 27160 11280
rect 26620 11240 27160 11268
rect 27154 11228 27160 11240
rect 27212 11268 27218 11280
rect 27433 11271 27491 11277
rect 27433 11268 27445 11271
rect 27212 11240 27445 11268
rect 27212 11228 27218 11240
rect 27433 11237 27445 11240
rect 27479 11237 27491 11271
rect 27433 11231 27491 11237
rect 27522 11228 27528 11280
rect 27580 11268 27586 11280
rect 28721 11271 28779 11277
rect 28721 11268 28733 11271
rect 27580 11240 28733 11268
rect 27580 11228 27586 11240
rect 28721 11237 28733 11240
rect 28767 11237 28779 11271
rect 28721 11231 28779 11237
rect 28810 11228 28816 11280
rect 28868 11268 28874 11280
rect 29825 11271 29883 11277
rect 29825 11268 29837 11271
rect 28868 11240 29837 11268
rect 28868 11228 28874 11240
rect 29825 11237 29837 11240
rect 29871 11237 29883 11271
rect 29825 11231 29883 11237
rect 32030 11228 32036 11280
rect 32088 11228 32094 11280
rect 32398 11228 32404 11280
rect 32456 11268 32462 11280
rect 32582 11268 32588 11280
rect 32456 11240 32588 11268
rect 32456 11228 32462 11240
rect 32582 11228 32588 11240
rect 32640 11228 32646 11280
rect 34146 11228 34152 11280
rect 34204 11268 34210 11280
rect 34333 11271 34391 11277
rect 34333 11268 34345 11271
rect 34204 11240 34345 11268
rect 34204 11228 34210 11240
rect 34333 11237 34345 11240
rect 34379 11268 34391 11271
rect 35986 11268 35992 11280
rect 34379 11240 35992 11268
rect 34379 11237 34391 11240
rect 34333 11231 34391 11237
rect 35986 11228 35992 11240
rect 36044 11228 36050 11280
rect 26602 11160 26608 11212
rect 26660 11200 26666 11212
rect 26660 11172 26740 11200
rect 26660 11160 26666 11172
rect 26712 11141 26740 11172
rect 27890 11160 27896 11212
rect 27948 11160 27954 11212
rect 27985 11203 28043 11209
rect 27985 11169 27997 11203
rect 28031 11200 28043 11203
rect 30374 11200 30380 11212
rect 28031 11172 30380 11200
rect 28031 11169 28043 11172
rect 27985 11163 28043 11169
rect 30374 11160 30380 11172
rect 30432 11160 30438 11212
rect 31202 11160 31208 11212
rect 31260 11160 31266 11212
rect 31389 11203 31447 11209
rect 31389 11169 31401 11203
rect 31435 11200 31447 11203
rect 31754 11200 31760 11212
rect 31435 11172 31760 11200
rect 31435 11169 31447 11172
rect 31389 11163 31447 11169
rect 31754 11160 31760 11172
rect 31812 11160 31818 11212
rect 31956 11172 34928 11200
rect 26375 11104 26464 11132
rect 26513 11135 26571 11141
rect 26375 11101 26387 11104
rect 26329 11095 26387 11101
rect 26513 11101 26525 11135
rect 26559 11101 26571 11135
rect 26513 11095 26571 11101
rect 26697 11135 26755 11141
rect 26697 11101 26709 11135
rect 26743 11101 26755 11135
rect 26697 11095 26755 11101
rect 26878 11092 26884 11144
rect 26936 11132 26942 11144
rect 28534 11132 28540 11144
rect 26936 11104 28540 11132
rect 26936 11092 26942 11104
rect 28534 11092 28540 11104
rect 28592 11092 28598 11144
rect 28629 11135 28687 11141
rect 28629 11101 28641 11135
rect 28675 11132 28687 11135
rect 28718 11132 28724 11144
rect 28675 11104 28724 11132
rect 28675 11101 28687 11104
rect 28629 11095 28687 11101
rect 28718 11092 28724 11104
rect 28776 11092 28782 11144
rect 29733 11135 29791 11141
rect 29733 11101 29745 11135
rect 29779 11132 29791 11135
rect 30006 11132 30012 11144
rect 29779 11104 30012 11132
rect 29779 11101 29791 11104
rect 29733 11095 29791 11101
rect 30006 11092 30012 11104
rect 30064 11132 30070 11144
rect 30190 11132 30196 11144
rect 30064 11104 30196 11132
rect 30064 11092 30070 11104
rect 30190 11092 30196 11104
rect 30248 11132 30254 11144
rect 31956 11141 31984 11172
rect 31941 11135 31999 11141
rect 31941 11132 31953 11135
rect 30248 11104 31953 11132
rect 30248 11092 30254 11104
rect 31941 11101 31953 11104
rect 31987 11101 31999 11135
rect 31941 11095 31999 11101
rect 32582 11092 32588 11144
rect 32640 11092 32646 11144
rect 34900 11141 34928 11172
rect 36262 11160 36268 11212
rect 36320 11200 36326 11212
rect 38565 11203 38623 11209
rect 38565 11200 38577 11203
rect 36320 11172 38577 11200
rect 36320 11160 36326 11172
rect 38565 11169 38577 11172
rect 38611 11169 38623 11203
rect 38565 11163 38623 11169
rect 34885 11135 34943 11141
rect 34885 11101 34897 11135
rect 34931 11101 34943 11135
rect 34885 11095 34943 11101
rect 35529 11135 35587 11141
rect 35529 11101 35541 11135
rect 35575 11132 35587 11135
rect 36173 11135 36231 11141
rect 36173 11132 36185 11135
rect 35575 11104 36185 11132
rect 35575 11101 35587 11104
rect 35529 11095 35587 11101
rect 36173 11101 36185 11104
rect 36219 11132 36231 11135
rect 36817 11135 36875 11141
rect 36817 11132 36829 11135
rect 36219 11104 36829 11132
rect 36219 11101 36231 11104
rect 36173 11095 36231 11101
rect 36817 11101 36829 11104
rect 36863 11132 36875 11135
rect 37458 11132 37464 11144
rect 36863 11104 37464 11132
rect 36863 11101 36875 11104
rect 36817 11095 36875 11101
rect 37458 11092 37464 11104
rect 37516 11132 37522 11144
rect 37553 11135 37611 11141
rect 37553 11132 37565 11135
rect 37516 11104 37565 11132
rect 37516 11092 37522 11104
rect 37553 11101 37565 11104
rect 37599 11132 37611 11135
rect 38102 11132 38108 11144
rect 37599 11104 38108 11132
rect 37599 11101 37611 11104
rect 37553 11095 37611 11101
rect 38102 11092 38108 11104
rect 38160 11092 38166 11144
rect 26418 11064 26424 11076
rect 24360 11036 24716 11064
rect 25148 11036 26424 11064
rect 24360 11024 24366 11036
rect 14568 10968 14780 10996
rect 16758 10956 16764 11008
rect 16816 10956 16822 11008
rect 17126 10956 17132 11008
rect 17184 10956 17190 11008
rect 19426 10956 19432 11008
rect 19484 10956 19490 11008
rect 19521 10999 19579 11005
rect 19521 10965 19533 10999
rect 19567 10996 19579 10999
rect 21726 10996 21732 11008
rect 19567 10968 21732 10996
rect 19567 10965 19579 10968
rect 19521 10959 19579 10965
rect 21726 10956 21732 10968
rect 21784 10956 21790 11008
rect 22097 10999 22155 11005
rect 22097 10965 22109 10999
rect 22143 10996 22155 10999
rect 24210 10996 24216 11008
rect 22143 10968 24216 10996
rect 22143 10965 22155 10968
rect 22097 10959 22155 10965
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 25148 11005 25176 11036
rect 26418 11024 26424 11036
rect 26476 11024 26482 11076
rect 26605 11067 26663 11073
rect 26605 11033 26617 11067
rect 26651 11033 26663 11067
rect 26605 11027 26663 11033
rect 25133 10999 25191 11005
rect 25133 10965 25145 10999
rect 25179 10965 25191 10999
rect 25133 10959 25191 10965
rect 25590 10956 25596 11008
rect 25648 10956 25654 11008
rect 25774 10956 25780 11008
rect 25832 10996 25838 11008
rect 26620 10996 26648 11027
rect 26786 11024 26792 11076
rect 26844 11064 26850 11076
rect 27433 11067 27491 11073
rect 27433 11064 27445 11067
rect 26844 11036 27445 11064
rect 26844 11024 26850 11036
rect 27433 11033 27445 11036
rect 27479 11064 27491 11067
rect 27706 11064 27712 11076
rect 27479 11036 27712 11064
rect 27479 11033 27491 11036
rect 27433 11027 27491 11033
rect 27706 11024 27712 11036
rect 27764 11024 27770 11076
rect 28552 11064 28580 11092
rect 29178 11064 29184 11076
rect 28092 11036 28304 11064
rect 28552 11036 29184 11064
rect 25832 10968 26648 10996
rect 25832 10956 25838 10968
rect 26878 10956 26884 11008
rect 26936 10956 26942 11008
rect 27154 10956 27160 11008
rect 27212 10996 27218 11008
rect 28092 10996 28120 11036
rect 27212 10968 28120 10996
rect 27212 10956 27218 10968
rect 28166 10956 28172 11008
rect 28224 10956 28230 11008
rect 28276 10996 28304 11036
rect 29178 11024 29184 11036
rect 29236 11024 29242 11076
rect 29638 11024 29644 11076
rect 29696 11064 29702 11076
rect 31018 11064 31024 11076
rect 29696 11036 31024 11064
rect 29696 11024 29702 11036
rect 31018 11024 31024 11036
rect 31076 11024 31082 11076
rect 31113 11067 31171 11073
rect 31113 11033 31125 11067
rect 31159 11064 31171 11067
rect 31294 11064 31300 11076
rect 31159 11036 31300 11064
rect 31159 11033 31171 11036
rect 31113 11027 31171 11033
rect 31294 11024 31300 11036
rect 31352 11064 31358 11076
rect 31570 11064 31576 11076
rect 31352 11036 31576 11064
rect 31352 11024 31358 11036
rect 31570 11024 31576 11036
rect 31628 11024 31634 11076
rect 32858 11024 32864 11076
rect 32916 11024 32922 11076
rect 33870 11024 33876 11076
rect 33928 11024 33934 11076
rect 34422 11024 34428 11076
rect 34480 11064 34486 11076
rect 35621 11067 35679 11073
rect 35621 11064 35633 11067
rect 34480 11036 35633 11064
rect 34480 11024 34486 11036
rect 35621 11033 35633 11036
rect 35667 11033 35679 11067
rect 35621 11027 35679 11033
rect 36372 11036 37044 11064
rect 30558 10996 30564 11008
rect 28276 10968 30564 10996
rect 30558 10956 30564 10968
rect 30616 10956 30622 11008
rect 31036 10996 31064 11024
rect 31478 10996 31484 11008
rect 31036 10968 31484 10996
rect 31478 10956 31484 10968
rect 31536 10956 31542 11008
rect 32122 10956 32128 11008
rect 32180 10996 32186 11008
rect 36372 10996 36400 11036
rect 32180 10968 36400 10996
rect 32180 10956 32186 10968
rect 36446 10956 36452 11008
rect 36504 10996 36510 11008
rect 36909 10999 36967 11005
rect 36909 10996 36921 10999
rect 36504 10968 36921 10996
rect 36504 10956 36510 10968
rect 36909 10965 36921 10968
rect 36955 10965 36967 10999
rect 37016 10996 37044 11036
rect 37642 11024 37648 11076
rect 37700 11024 37706 11076
rect 38289 11067 38347 11073
rect 38289 11033 38301 11067
rect 38335 11064 38347 11067
rect 39390 11064 39396 11076
rect 38335 11036 39396 11064
rect 38335 11033 38347 11036
rect 38289 11027 38347 11033
rect 39390 11024 39396 11036
rect 39448 11024 39454 11076
rect 37734 10996 37740 11008
rect 37016 10968 37740 10996
rect 36909 10959 36967 10965
rect 37734 10956 37740 10968
rect 37792 10956 37798 11008
rect 1104 10906 39352 10928
rect 1104 10854 10472 10906
rect 10524 10854 10536 10906
rect 10588 10854 10600 10906
rect 10652 10854 10664 10906
rect 10716 10854 10728 10906
rect 10780 10854 19994 10906
rect 20046 10854 20058 10906
rect 20110 10854 20122 10906
rect 20174 10854 20186 10906
rect 20238 10854 20250 10906
rect 20302 10854 29516 10906
rect 29568 10854 29580 10906
rect 29632 10854 29644 10906
rect 29696 10854 29708 10906
rect 29760 10854 29772 10906
rect 29824 10854 39038 10906
rect 39090 10854 39102 10906
rect 39154 10854 39166 10906
rect 39218 10854 39230 10906
rect 39282 10854 39294 10906
rect 39346 10854 39352 10906
rect 1104 10832 39352 10854
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 5258 10792 5264 10804
rect 2179 10764 5264 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5350 10752 5356 10804
rect 5408 10792 5414 10804
rect 5829 10795 5887 10801
rect 5829 10792 5841 10795
rect 5408 10764 5841 10792
rect 5408 10752 5414 10764
rect 5829 10761 5841 10764
rect 5875 10792 5887 10795
rect 7025 10795 7083 10801
rect 7025 10792 7037 10795
rect 5875 10764 7037 10792
rect 5875 10761 5887 10764
rect 5829 10755 5887 10761
rect 7025 10761 7037 10764
rect 7071 10792 7083 10795
rect 8202 10792 8208 10804
rect 7071 10764 8208 10792
rect 7071 10761 7083 10764
rect 7025 10755 7083 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 8904 10764 9352 10792
rect 8904 10752 8910 10764
rect 1946 10684 1952 10736
rect 2004 10724 2010 10736
rect 2041 10727 2099 10733
rect 2041 10724 2053 10727
rect 2004 10696 2053 10724
rect 2004 10684 2010 10696
rect 2041 10693 2053 10696
rect 2087 10693 2099 10727
rect 2041 10687 2099 10693
rect 2406 10684 2412 10736
rect 2464 10724 2470 10736
rect 5629 10727 5687 10733
rect 2464 10696 3634 10724
rect 2464 10684 2470 10696
rect 5629 10693 5641 10727
rect 5675 10724 5687 10727
rect 5718 10724 5724 10736
rect 5675 10696 5724 10724
rect 5675 10693 5687 10696
rect 5629 10687 5687 10693
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 6730 10684 6736 10736
rect 6788 10724 6794 10736
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 6788 10696 6837 10724
rect 6788 10684 6794 10696
rect 6825 10693 6837 10696
rect 6871 10693 6883 10727
rect 6825 10687 6883 10693
rect 7929 10727 7987 10733
rect 7929 10693 7941 10727
rect 7975 10724 7987 10727
rect 8018 10724 8024 10736
rect 7975 10696 8024 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 9324 10724 9352 10764
rect 9398 10752 9404 10804
rect 9456 10792 9462 10804
rect 9456 10764 10548 10792
rect 9456 10752 9462 10764
rect 9677 10727 9735 10733
rect 9677 10724 9689 10727
rect 9324 10696 9689 10724
rect 9677 10693 9689 10696
rect 9723 10693 9735 10727
rect 9677 10687 9735 10693
rect 10042 10684 10048 10736
rect 10100 10724 10106 10736
rect 10413 10727 10471 10733
rect 10413 10724 10425 10727
rect 10100 10696 10425 10724
rect 10100 10684 10106 10696
rect 10413 10693 10425 10696
rect 10459 10693 10471 10727
rect 10413 10687 10471 10693
rect 2866 10616 2872 10668
rect 2924 10616 2930 10668
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7650 10656 7656 10668
rect 6972 10628 7656 10656
rect 6972 10616 6978 10628
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 9030 10616 9036 10668
rect 9088 10616 9094 10668
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 10137 10659 10195 10665
rect 10137 10656 10149 10659
rect 9456 10628 10149 10656
rect 9456 10616 9462 10628
rect 10137 10625 10149 10628
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10520 10665 10548 10764
rect 11900 10764 14412 10792
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 10284 10628 10333 10656
rect 10284 10616 10290 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 11054 10656 11060 10668
rect 10551 10628 11060 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11698 10616 11704 10668
rect 11756 10616 11762 10668
rect 11900 10665 11928 10764
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12989 10727 13047 10733
rect 12989 10724 13001 10727
rect 12124 10696 13001 10724
rect 12124 10684 12130 10696
rect 12989 10693 13001 10696
rect 13035 10693 13047 10727
rect 12989 10687 13047 10693
rect 13446 10684 13452 10736
rect 13504 10684 13510 10736
rect 14384 10724 14412 10764
rect 14458 10752 14464 10804
rect 14516 10752 14522 10804
rect 14918 10752 14924 10804
rect 14976 10792 14982 10804
rect 15378 10792 15384 10804
rect 14976 10764 15384 10792
rect 14976 10752 14982 10764
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 17221 10795 17279 10801
rect 15620 10764 16804 10792
rect 15620 10752 15626 10764
rect 16666 10724 16672 10736
rect 14384 10696 16672 10724
rect 16666 10684 16672 10696
rect 16724 10684 16730 10736
rect 16776 10724 16804 10764
rect 17221 10761 17233 10795
rect 17267 10761 17279 10795
rect 17221 10755 17279 10761
rect 17313 10795 17371 10801
rect 17313 10761 17325 10795
rect 17359 10792 17371 10795
rect 18598 10792 18604 10804
rect 17359 10764 18604 10792
rect 17359 10761 17371 10764
rect 17313 10755 17371 10761
rect 17236 10724 17264 10755
rect 18598 10752 18604 10764
rect 18656 10792 18662 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 18656 10764 19809 10792
rect 18656 10752 18662 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 22097 10795 22155 10801
rect 22097 10761 22109 10795
rect 22143 10792 22155 10795
rect 22278 10792 22284 10804
rect 22143 10764 22284 10792
rect 22143 10761 22155 10764
rect 22097 10755 22155 10761
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 23842 10792 23848 10804
rect 22664 10764 23848 10792
rect 16776 10696 17264 10724
rect 17494 10684 17500 10736
rect 17552 10724 17558 10736
rect 18325 10727 18383 10733
rect 18325 10724 18337 10727
rect 17552 10696 18337 10724
rect 17552 10684 17558 10696
rect 18325 10693 18337 10696
rect 18371 10693 18383 10727
rect 21358 10724 21364 10736
rect 19550 10696 21364 10724
rect 18325 10687 18383 10693
rect 21358 10684 21364 10696
rect 21416 10684 21422 10736
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10656 15531 10659
rect 15519 10628 17816 10656
rect 15519 10625 15531 10628
rect 15473 10619 15531 10625
rect 2314 10548 2320 10600
rect 2372 10588 2378 10600
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 2372 10560 3157 10588
rect 2372 10548 2378 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 3145 10551 3203 10557
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 12618 10588 12624 10600
rect 3936 10560 5856 10588
rect 3936 10548 3942 10560
rect 3786 10412 3792 10464
rect 3844 10452 3850 10464
rect 5828 10461 5856 10560
rect 9048 10560 12624 10588
rect 5994 10480 6000 10532
rect 6052 10480 6058 10532
rect 8938 10480 8944 10532
rect 8996 10520 9002 10532
rect 9048 10520 9076 10560
rect 12618 10548 12624 10560
rect 12676 10548 12682 10600
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 8996 10492 9076 10520
rect 8996 10480 9002 10492
rect 9122 10480 9128 10532
rect 9180 10520 9186 10532
rect 10226 10520 10232 10532
rect 9180 10492 10232 10520
rect 9180 10480 9186 10492
rect 10226 10480 10232 10492
rect 10284 10480 10290 10532
rect 10612 10492 11744 10520
rect 4617 10455 4675 10461
rect 4617 10452 4629 10455
rect 3844 10424 4629 10452
rect 3844 10412 3850 10424
rect 4617 10421 4629 10424
rect 4663 10421 4675 10455
rect 4617 10415 4675 10421
rect 5813 10455 5871 10461
rect 5813 10421 5825 10455
rect 5859 10452 5871 10455
rect 7009 10455 7067 10461
rect 7009 10452 7021 10455
rect 5859 10424 7021 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 7009 10421 7021 10424
rect 7055 10452 7067 10455
rect 7098 10452 7104 10464
rect 7055 10424 7104 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7193 10455 7251 10461
rect 7193 10421 7205 10455
rect 7239 10452 7251 10455
rect 10612 10452 10640 10492
rect 7239 10424 10640 10452
rect 10689 10455 10747 10461
rect 7239 10421 7251 10424
rect 7193 10415 7251 10421
rect 10689 10421 10701 10455
rect 10735 10452 10747 10455
rect 11422 10452 11428 10464
rect 10735 10424 11428 10452
rect 10735 10421 10747 10424
rect 10689 10415 10747 10421
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 11716 10461 11744 10492
rect 11701 10455 11759 10461
rect 11701 10421 11713 10455
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 12066 10412 12072 10464
rect 12124 10412 12130 10464
rect 12728 10452 12756 10551
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 13504 10560 14044 10588
rect 13504 10548 13510 10560
rect 14016 10520 14044 10560
rect 14458 10548 14464 10600
rect 14516 10588 14522 10600
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 14516 10560 15577 10588
rect 14516 10548 14522 10560
rect 15565 10557 15577 10560
rect 15611 10588 15623 10591
rect 16482 10588 16488 10600
rect 15611 10560 16488 10588
rect 15611 10557 15623 10560
rect 15565 10551 15623 10557
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 17310 10588 17316 10600
rect 16592 10560 17316 10588
rect 16592 10520 16620 10560
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 17402 10548 17408 10600
rect 17460 10548 17466 10600
rect 14016 10492 16620 10520
rect 16853 10523 16911 10529
rect 16853 10489 16865 10523
rect 16899 10520 16911 10523
rect 17494 10520 17500 10532
rect 16899 10492 17500 10520
rect 16899 10489 16911 10492
rect 16853 10483 16911 10489
rect 17494 10480 17500 10492
rect 17552 10480 17558 10532
rect 13722 10452 13728 10464
rect 12728 10424 13728 10452
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 15013 10455 15071 10461
rect 15013 10421 15025 10455
rect 15059 10452 15071 10455
rect 17126 10452 17132 10464
rect 15059 10424 17132 10452
rect 15059 10421 15071 10424
rect 15013 10415 15071 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17788 10452 17816 10628
rect 19794 10616 19800 10668
rect 19852 10656 19858 10668
rect 20349 10659 20407 10665
rect 20349 10656 20361 10659
rect 19852 10628 20361 10656
rect 19852 10616 19858 10628
rect 20349 10625 20361 10628
rect 20395 10625 20407 10659
rect 20349 10619 20407 10625
rect 20622 10616 20628 10668
rect 20680 10656 20686 10668
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 20680 10628 22017 10656
rect 20680 10616 20686 10628
rect 22005 10625 22017 10628
rect 22051 10656 22063 10659
rect 22664 10656 22692 10764
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 23934 10752 23940 10804
rect 23992 10792 23998 10804
rect 25501 10795 25559 10801
rect 25501 10792 25513 10795
rect 23992 10764 25513 10792
rect 23992 10752 23998 10764
rect 25501 10761 25513 10764
rect 25547 10761 25559 10795
rect 25958 10792 25964 10804
rect 25501 10755 25559 10761
rect 25608 10764 25964 10792
rect 24762 10724 24768 10736
rect 24150 10696 24768 10724
rect 24762 10684 24768 10696
rect 24820 10684 24826 10736
rect 25133 10727 25191 10733
rect 25133 10693 25145 10727
rect 25179 10693 25191 10727
rect 25133 10690 25191 10693
rect 25333 10727 25391 10733
rect 25333 10693 25345 10727
rect 25379 10724 25391 10727
rect 25608 10724 25636 10764
rect 25958 10752 25964 10764
rect 26016 10752 26022 10804
rect 27157 10795 27215 10801
rect 27157 10761 27169 10795
rect 27203 10792 27215 10795
rect 27203 10764 28948 10792
rect 27203 10761 27215 10764
rect 27157 10755 27215 10761
rect 28166 10724 28172 10736
rect 25379 10696 25636 10724
rect 25992 10696 28172 10724
rect 25379 10693 25391 10696
rect 25133 10687 25202 10690
rect 25333 10687 25391 10693
rect 25148 10662 25202 10687
rect 22051 10628 22692 10656
rect 25174 10656 25202 10662
rect 25590 10656 25596 10668
rect 25174 10628 25596 10656
rect 22051 10625 22063 10628
rect 22005 10619 22063 10625
rect 25590 10616 25596 10628
rect 25648 10616 25654 10668
rect 25992 10665 26020 10696
rect 28166 10684 28172 10696
rect 28224 10684 28230 10736
rect 28920 10724 28948 10764
rect 29270 10752 29276 10804
rect 29328 10792 29334 10804
rect 30561 10795 30619 10801
rect 30561 10792 30573 10795
rect 29328 10764 30573 10792
rect 29328 10752 29334 10764
rect 30561 10761 30573 10764
rect 30607 10761 30619 10795
rect 30561 10755 30619 10761
rect 31021 10795 31079 10801
rect 31021 10761 31033 10795
rect 31067 10792 31079 10795
rect 32674 10792 32680 10804
rect 31067 10764 32680 10792
rect 31067 10761 31079 10764
rect 31021 10755 31079 10761
rect 32674 10752 32680 10764
rect 32732 10752 32738 10804
rect 33594 10752 33600 10804
rect 33652 10792 33658 10804
rect 33870 10792 33876 10804
rect 33652 10764 33876 10792
rect 33652 10752 33658 10764
rect 33870 10752 33876 10764
rect 33928 10752 33934 10804
rect 34974 10752 34980 10804
rect 35032 10792 35038 10804
rect 35710 10792 35716 10804
rect 35032 10764 35716 10792
rect 35032 10752 35038 10764
rect 35710 10752 35716 10764
rect 35768 10752 35774 10804
rect 29089 10727 29147 10733
rect 29089 10724 29101 10727
rect 28920 10696 29101 10724
rect 29089 10693 29101 10696
rect 29135 10693 29147 10727
rect 29089 10687 29147 10693
rect 29546 10684 29552 10736
rect 29604 10684 29610 10736
rect 32306 10684 32312 10736
rect 32364 10724 32370 10736
rect 32585 10727 32643 10733
rect 32585 10724 32597 10727
rect 32364 10696 32597 10724
rect 32364 10684 32370 10696
rect 32585 10693 32597 10696
rect 32631 10693 32643 10727
rect 34422 10724 34428 10736
rect 33810 10696 34428 10724
rect 32585 10687 32643 10693
rect 34422 10684 34428 10696
rect 34480 10684 34486 10736
rect 37366 10724 37372 10736
rect 36018 10696 37372 10724
rect 37366 10684 37372 10696
rect 37424 10684 37430 10736
rect 25961 10659 26020 10665
rect 25961 10625 25973 10659
rect 26007 10626 26020 10659
rect 26054 10659 26112 10665
rect 26007 10625 26019 10626
rect 25961 10619 26019 10625
rect 26054 10625 26066 10659
rect 26100 10625 26112 10659
rect 26054 10619 26112 10625
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17920 10560 18061 10588
rect 17920 10548 17926 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 20901 10591 20959 10597
rect 20901 10557 20913 10591
rect 20947 10588 20959 10591
rect 21266 10588 21272 10600
rect 20947 10560 21272 10588
rect 20947 10557 20959 10560
rect 20901 10551 20959 10557
rect 21266 10548 21272 10560
rect 21324 10548 21330 10600
rect 22649 10591 22707 10597
rect 22649 10557 22661 10591
rect 22695 10557 22707 10591
rect 22649 10551 22707 10557
rect 22925 10591 22983 10597
rect 22925 10557 22937 10591
rect 22971 10588 22983 10591
rect 24486 10588 24492 10600
rect 22971 10560 24492 10588
rect 22971 10557 22983 10560
rect 22925 10551 22983 10557
rect 20622 10480 20628 10532
rect 20680 10520 20686 10532
rect 22664 10520 22692 10551
rect 24486 10548 24492 10560
rect 24544 10548 24550 10600
rect 24673 10591 24731 10597
rect 24673 10557 24685 10591
rect 24719 10588 24731 10591
rect 25038 10588 25044 10600
rect 24719 10560 25044 10588
rect 24719 10557 24731 10560
rect 24673 10551 24731 10557
rect 25038 10548 25044 10560
rect 25096 10548 25102 10600
rect 25130 10548 25136 10600
rect 25188 10588 25194 10600
rect 26069 10588 26097 10619
rect 26234 10616 26240 10668
rect 26292 10616 26298 10668
rect 26326 10616 26332 10668
rect 26384 10616 26390 10668
rect 26467 10659 26525 10665
rect 26467 10625 26479 10659
rect 26513 10656 26525 10659
rect 27062 10656 27068 10668
rect 26513 10628 27068 10656
rect 26513 10625 26525 10628
rect 26467 10619 26525 10625
rect 27062 10616 27068 10628
rect 27120 10616 27126 10668
rect 27430 10616 27436 10668
rect 27488 10656 27494 10668
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 27488 10628 27537 10656
rect 27488 10616 27494 10628
rect 27525 10625 27537 10628
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 27617 10659 27675 10665
rect 27617 10625 27629 10659
rect 27663 10656 27675 10659
rect 28258 10656 28264 10668
rect 27663 10628 28264 10656
rect 27663 10625 27675 10628
rect 27617 10619 27675 10625
rect 28258 10616 28264 10628
rect 28316 10616 28322 10668
rect 30558 10616 30564 10668
rect 30616 10656 30622 10668
rect 31386 10656 31392 10668
rect 30616 10628 31392 10656
rect 30616 10616 30622 10628
rect 31386 10616 31392 10628
rect 31444 10616 31450 10668
rect 31846 10656 31852 10668
rect 31496 10628 31852 10656
rect 26694 10588 26700 10600
rect 25188 10560 26097 10588
rect 26528 10560 26700 10588
rect 25188 10548 25194 10560
rect 20680 10492 22692 10520
rect 20680 10480 20686 10492
rect 18782 10452 18788 10464
rect 17788 10424 18788 10452
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 22664 10452 22692 10492
rect 24394 10480 24400 10532
rect 24452 10520 24458 10532
rect 26528 10520 26556 10560
rect 26694 10548 26700 10560
rect 26752 10588 26758 10600
rect 27246 10588 27252 10600
rect 26752 10560 27252 10588
rect 26752 10548 26758 10560
rect 27246 10548 27252 10560
rect 27304 10588 27310 10600
rect 27709 10591 27767 10597
rect 27709 10588 27721 10591
rect 27304 10560 27721 10588
rect 27304 10548 27310 10560
rect 27709 10557 27721 10560
rect 27755 10557 27767 10591
rect 27709 10551 27767 10557
rect 28813 10591 28871 10597
rect 28813 10557 28825 10591
rect 28859 10557 28871 10591
rect 28813 10551 28871 10557
rect 24452 10492 26556 10520
rect 26605 10523 26663 10529
rect 24452 10480 24458 10492
rect 26605 10489 26617 10523
rect 26651 10520 26663 10523
rect 27154 10520 27160 10532
rect 26651 10492 27160 10520
rect 26651 10489 26663 10492
rect 26605 10483 26663 10489
rect 27154 10480 27160 10492
rect 27212 10480 27218 10532
rect 23658 10452 23664 10464
rect 22664 10424 23664 10452
rect 23658 10412 23664 10424
rect 23716 10412 23722 10464
rect 25317 10455 25375 10461
rect 25317 10421 25329 10455
rect 25363 10452 25375 10455
rect 25498 10452 25504 10464
rect 25363 10424 25504 10452
rect 25363 10421 25375 10424
rect 25317 10415 25375 10421
rect 25498 10412 25504 10424
rect 25556 10412 25562 10464
rect 25590 10412 25596 10464
rect 25648 10452 25654 10464
rect 26234 10452 26240 10464
rect 25648 10424 26240 10452
rect 25648 10412 25654 10424
rect 26234 10412 26240 10424
rect 26292 10452 26298 10464
rect 28074 10452 28080 10464
rect 26292 10424 28080 10452
rect 26292 10412 26298 10424
rect 28074 10412 28080 10424
rect 28132 10412 28138 10464
rect 28828 10452 28856 10551
rect 29086 10548 29092 10600
rect 29144 10588 29150 10600
rect 31496 10597 31524 10628
rect 31846 10616 31852 10628
rect 31904 10616 31910 10668
rect 34514 10616 34520 10668
rect 34572 10616 34578 10668
rect 36725 10659 36783 10665
rect 36725 10625 36737 10659
rect 36771 10656 36783 10659
rect 37461 10659 37519 10665
rect 37461 10656 37473 10659
rect 36771 10628 37473 10656
rect 36771 10625 36783 10628
rect 36725 10619 36783 10625
rect 37461 10625 37473 10628
rect 37507 10656 37519 10659
rect 37826 10656 37832 10668
rect 37507 10628 37832 10656
rect 37507 10625 37519 10628
rect 37461 10619 37519 10625
rect 37826 10616 37832 10628
rect 37884 10656 37890 10668
rect 38010 10656 38016 10668
rect 37884 10628 38016 10656
rect 37884 10616 37890 10628
rect 38010 10616 38016 10628
rect 38068 10616 38074 10668
rect 38105 10659 38163 10665
rect 38105 10625 38117 10659
rect 38151 10656 38163 10659
rect 38378 10656 38384 10668
rect 38151 10628 38384 10656
rect 38151 10625 38163 10628
rect 38105 10619 38163 10625
rect 38378 10616 38384 10628
rect 38436 10616 38442 10668
rect 31481 10591 31539 10597
rect 31481 10588 31493 10591
rect 29144 10560 31493 10588
rect 29144 10548 29150 10560
rect 31481 10557 31493 10560
rect 31527 10557 31539 10591
rect 31481 10551 31539 10557
rect 31573 10591 31631 10597
rect 31573 10557 31585 10591
rect 31619 10557 31631 10591
rect 31573 10551 31631 10557
rect 32309 10591 32367 10597
rect 32309 10557 32321 10591
rect 32355 10588 32367 10591
rect 32582 10588 32588 10600
rect 32355 10560 32588 10588
rect 32355 10557 32367 10560
rect 32309 10551 32367 10557
rect 30466 10480 30472 10532
rect 30524 10520 30530 10532
rect 31202 10520 31208 10532
rect 30524 10492 31208 10520
rect 30524 10480 30530 10492
rect 31202 10480 31208 10492
rect 31260 10520 31266 10532
rect 31588 10520 31616 10551
rect 32582 10548 32588 10560
rect 32640 10548 32646 10600
rect 34790 10548 34796 10600
rect 34848 10548 34854 10600
rect 31260 10492 31616 10520
rect 31260 10480 31266 10492
rect 33686 10480 33692 10532
rect 33744 10520 33750 10532
rect 34146 10520 34152 10532
rect 33744 10492 34152 10520
rect 33744 10480 33750 10492
rect 34146 10480 34152 10492
rect 34204 10480 34210 10532
rect 30190 10452 30196 10464
rect 28828 10424 30196 10452
rect 30190 10412 30196 10424
rect 30248 10412 30254 10464
rect 31386 10412 31392 10464
rect 31444 10452 31450 10464
rect 32122 10452 32128 10464
rect 31444 10424 32128 10452
rect 31444 10412 31450 10424
rect 32122 10412 32128 10424
rect 32180 10412 32186 10464
rect 33594 10412 33600 10464
rect 33652 10452 33658 10464
rect 34057 10455 34115 10461
rect 34057 10452 34069 10455
rect 33652 10424 34069 10452
rect 33652 10412 33658 10424
rect 34057 10421 34069 10424
rect 34103 10421 34115 10455
rect 34057 10415 34115 10421
rect 35802 10412 35808 10464
rect 35860 10452 35866 10464
rect 36265 10455 36323 10461
rect 36265 10452 36277 10455
rect 35860 10424 36277 10452
rect 35860 10412 35866 10424
rect 36265 10421 36277 10424
rect 36311 10421 36323 10455
rect 36265 10415 36323 10421
rect 36630 10412 36636 10464
rect 36688 10452 36694 10464
rect 36817 10455 36875 10461
rect 36817 10452 36829 10455
rect 36688 10424 36829 10452
rect 36688 10412 36694 10424
rect 36817 10421 36829 10424
rect 36863 10421 36875 10455
rect 36817 10415 36875 10421
rect 37553 10455 37611 10461
rect 37553 10421 37565 10455
rect 37599 10452 37611 10455
rect 37642 10452 37648 10464
rect 37599 10424 37648 10452
rect 37599 10421 37611 10424
rect 37553 10415 37611 10421
rect 37642 10412 37648 10424
rect 37700 10412 37706 10464
rect 38194 10412 38200 10464
rect 38252 10412 38258 10464
rect 1104 10362 39192 10384
rect 1104 10310 5711 10362
rect 5763 10310 5775 10362
rect 5827 10310 5839 10362
rect 5891 10310 5903 10362
rect 5955 10310 5967 10362
rect 6019 10310 15233 10362
rect 15285 10310 15297 10362
rect 15349 10310 15361 10362
rect 15413 10310 15425 10362
rect 15477 10310 15489 10362
rect 15541 10310 24755 10362
rect 24807 10310 24819 10362
rect 24871 10310 24883 10362
rect 24935 10310 24947 10362
rect 24999 10310 25011 10362
rect 25063 10310 34277 10362
rect 34329 10310 34341 10362
rect 34393 10310 34405 10362
rect 34457 10310 34469 10362
rect 34521 10310 34533 10362
rect 34585 10310 39192 10362
rect 1104 10288 39192 10310
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 5350 10248 5356 10260
rect 2740 10220 5356 10248
rect 2740 10208 2746 10220
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 5626 10208 5632 10260
rect 5684 10208 5690 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 8938 10248 8944 10260
rect 8619 10220 8944 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 10042 10248 10048 10260
rect 9732 10220 10048 10248
rect 9732 10208 9738 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 12529 10251 12587 10257
rect 12529 10248 12541 10251
rect 10284 10220 12541 10248
rect 10284 10208 10290 10220
rect 12529 10217 12541 10220
rect 12575 10217 12587 10251
rect 14090 10248 14096 10260
rect 12529 10211 12587 10217
rect 12728 10220 14096 10248
rect 9306 10180 9312 10192
rect 8128 10152 9312 10180
rect 2590 10112 2596 10124
rect 2332 10084 2596 10112
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 2332 10053 2360 10084
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 4890 10112 4896 10124
rect 4847 10084 4896 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 6546 10112 6552 10124
rect 5868 10084 6552 10112
rect 5868 10072 5874 10084
rect 6546 10072 6552 10084
rect 6604 10112 6610 10124
rect 8128 10112 8156 10152
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 11054 10140 11060 10192
rect 11112 10180 11118 10192
rect 12728 10180 12756 10220
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 14366 10208 14372 10260
rect 14424 10208 14430 10260
rect 15013 10251 15071 10257
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 15059 10220 18092 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 11112 10152 12756 10180
rect 11112 10140 11118 10152
rect 6604 10084 8156 10112
rect 6604 10072 6610 10084
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 8904 10084 12296 10112
rect 8904 10072 8910 10084
rect 2317 10047 2375 10053
rect 2317 10044 2329 10047
rect 1820 10016 2329 10044
rect 1820 10004 1826 10016
rect 2317 10013 2329 10016
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 5166 10044 5172 10056
rect 3467 10016 5172 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5592 10016 6193 10044
rect 5592 10004 5598 10016
rect 6181 10013 6193 10016
rect 6227 10044 6239 10047
rect 6270 10044 6276 10056
rect 6227 10016 6276 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 6822 10004 6828 10056
rect 6880 10004 6886 10056
rect 8202 10004 8208 10056
rect 8260 10004 8266 10056
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 9585 10047 9643 10053
rect 9585 10044 9597 10047
rect 9364 10016 9597 10044
rect 9364 10004 9370 10016
rect 9585 10013 9597 10016
rect 9631 10013 9643 10047
rect 9585 10007 9643 10013
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 12268 10053 12296 10084
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 11388 10016 11989 10044
rect 11388 10004 11394 10016
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10044 12403 10047
rect 12728 10044 12756 10152
rect 12894 10140 12900 10192
rect 12952 10180 12958 10192
rect 12989 10183 13047 10189
rect 12989 10180 13001 10183
rect 12952 10152 13001 10180
rect 12952 10140 12958 10152
rect 12989 10149 13001 10152
rect 13035 10149 13047 10183
rect 12989 10143 13047 10149
rect 13078 10140 13084 10192
rect 13136 10180 13142 10192
rect 16482 10180 16488 10192
rect 13136 10152 16488 10180
rect 13136 10140 13142 10152
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 13648 10121 13676 10152
rect 16482 10140 16488 10152
rect 16540 10140 16546 10192
rect 16758 10140 16764 10192
rect 16816 10140 16822 10192
rect 18064 10180 18092 10220
rect 18506 10208 18512 10260
rect 18564 10208 18570 10260
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 26973 10251 27031 10257
rect 26973 10248 26985 10251
rect 20772 10220 26985 10248
rect 20772 10208 20778 10220
rect 26973 10217 26985 10220
rect 27019 10217 27031 10251
rect 30377 10251 30435 10257
rect 30377 10248 30389 10251
rect 26973 10211 27031 10217
rect 27080 10220 30389 10248
rect 18064 10152 20760 10180
rect 13449 10115 13507 10121
rect 13449 10112 13461 10115
rect 12860 10084 13461 10112
rect 12860 10072 12866 10084
rect 13449 10081 13461 10084
rect 13495 10081 13507 10115
rect 13449 10075 13507 10081
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10081 13691 10115
rect 14918 10112 14924 10124
rect 13633 10075 13691 10081
rect 14200 10084 14924 10112
rect 12391 10016 12756 10044
rect 13357 10047 13415 10053
rect 12391 10013 12403 10016
rect 12345 10007 12403 10013
rect 13357 10013 13369 10047
rect 13403 10044 13415 10047
rect 14200 10044 14228 10084
rect 14918 10072 14924 10084
rect 14976 10072 14982 10124
rect 15565 10115 15623 10121
rect 15565 10112 15577 10115
rect 15028 10084 15577 10112
rect 13403 10016 14228 10044
rect 14277 10047 14335 10053
rect 13403 10013 13415 10016
rect 13357 10007 13415 10013
rect 14277 10013 14289 10047
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 2222 9976 2228 9988
rect 1719 9948 2228 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 2222 9936 2228 9948
rect 2280 9936 2286 9988
rect 2590 9936 2596 9988
rect 2648 9936 2654 9988
rect 3237 9979 3295 9985
rect 3237 9945 3249 9979
rect 3283 9976 3295 9979
rect 4430 9976 4436 9988
rect 3283 9948 4436 9976
rect 3283 9945 3295 9948
rect 3237 9939 3295 9945
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 4617 9979 4675 9985
rect 4617 9945 4629 9979
rect 4663 9976 4675 9979
rect 6086 9976 6092 9988
rect 4663 9948 6092 9976
rect 4663 9945 4675 9948
rect 4617 9939 4675 9945
rect 6086 9936 6092 9948
rect 6144 9976 6150 9988
rect 6144 9948 6960 9976
rect 6144 9936 6150 9948
rect 6932 9920 6960 9948
rect 7098 9936 7104 9988
rect 7156 9936 7162 9988
rect 9858 9936 9864 9988
rect 9916 9936 9922 9988
rect 11146 9976 11152 9988
rect 11086 9948 11152 9976
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 11882 9936 11888 9988
rect 11940 9976 11946 9988
rect 12161 9979 12219 9985
rect 12161 9976 12173 9979
rect 11940 9948 12173 9976
rect 11940 9936 11946 9948
rect 12161 9945 12173 9948
rect 12207 9976 12219 9979
rect 13446 9976 13452 9988
rect 12207 9948 13452 9976
rect 12207 9945 12219 9948
rect 12161 9939 12219 9945
rect 13446 9936 13452 9948
rect 13504 9936 13510 9988
rect 13538 9936 13544 9988
rect 13596 9976 13602 9988
rect 14292 9976 14320 10007
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 15028 10044 15056 10084
rect 15565 10081 15577 10084
rect 15611 10081 15623 10115
rect 16776 10112 16804 10140
rect 17037 10115 17095 10121
rect 17037 10112 17049 10115
rect 16776 10084 17049 10112
rect 15565 10075 15623 10081
rect 17037 10081 17049 10084
rect 17083 10081 17095 10115
rect 17037 10075 17095 10081
rect 17402 10072 17408 10124
rect 17460 10112 17466 10124
rect 17678 10112 17684 10124
rect 17460 10084 17684 10112
rect 17460 10072 17466 10084
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 19702 10072 19708 10124
rect 19760 10112 19766 10124
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 19760 10084 19809 10112
rect 19760 10072 19766 10084
rect 19797 10081 19809 10084
rect 19843 10081 19855 10115
rect 19797 10075 19855 10081
rect 20622 10072 20628 10124
rect 20680 10072 20686 10124
rect 20732 10112 20760 10152
rect 24688 10152 24900 10180
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20732 10084 20913 10112
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 20901 10075 20959 10081
rect 21634 10072 21640 10124
rect 21692 10112 21698 10124
rect 21692 10084 22232 10112
rect 21692 10072 21698 10084
rect 16298 10044 16304 10056
rect 14884 10016 15056 10044
rect 15304 10016 16304 10044
rect 14884 10004 14890 10016
rect 15304 9976 15332 10016
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 16758 10004 16764 10056
rect 16816 10004 16822 10056
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19521 10047 19579 10053
rect 19521 10044 19533 10047
rect 19392 10016 19533 10044
rect 19392 10004 19398 10016
rect 19521 10013 19533 10016
rect 19567 10013 19579 10047
rect 19521 10007 19579 10013
rect 13596 9948 15332 9976
rect 15381 9979 15439 9985
rect 13596 9936 13602 9948
rect 15381 9945 15393 9979
rect 15427 9976 15439 9979
rect 15654 9976 15660 9988
rect 15427 9948 15660 9976
rect 15427 9945 15439 9948
rect 15381 9939 15439 9945
rect 15654 9936 15660 9948
rect 15712 9936 15718 9988
rect 16206 9936 16212 9988
rect 16264 9976 16270 9988
rect 16264 9948 17526 9976
rect 19812 9948 20852 9976
rect 16264 9936 16270 9948
rect 1026 9868 1032 9920
rect 1084 9908 1090 9920
rect 1765 9911 1823 9917
rect 1765 9908 1777 9911
rect 1084 9880 1777 9908
rect 1084 9868 1090 9880
rect 1765 9877 1777 9880
rect 1811 9877 1823 9911
rect 1765 9871 1823 9877
rect 4154 9868 4160 9920
rect 4212 9868 4218 9920
rect 4522 9868 4528 9920
rect 4580 9868 4586 9920
rect 6273 9911 6331 9917
rect 6273 9877 6285 9911
rect 6319 9908 6331 9911
rect 6638 9908 6644 9920
rect 6319 9880 6644 9908
rect 6319 9877 6331 9880
rect 6273 9871 6331 9877
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 6914 9868 6920 9920
rect 6972 9868 6978 9920
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 7834 9908 7840 9920
rect 7248 9880 7840 9908
rect 7248 9868 7254 9880
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8018 9868 8024 9920
rect 8076 9908 8082 9920
rect 9030 9908 9036 9920
rect 8076 9880 9036 9908
rect 8076 9868 8082 9880
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 11164 9908 11192 9936
rect 9355 9880 11192 9908
rect 11333 9911 11391 9917
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 11333 9877 11345 9911
rect 11379 9908 11391 9911
rect 12526 9908 12532 9920
rect 11379 9880 12532 9908
rect 11379 9877 11391 9880
rect 11333 9871 11391 9877
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 13906 9908 13912 9920
rect 12952 9880 13912 9908
rect 12952 9868 12958 9880
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 15473 9911 15531 9917
rect 15473 9877 15485 9911
rect 15519 9908 15531 9911
rect 16022 9908 16028 9920
rect 15519 9880 16028 9908
rect 15519 9877 15531 9880
rect 15473 9871 15531 9877
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 19812 9908 19840 9948
rect 17276 9880 19840 9908
rect 17276 9868 17282 9880
rect 19886 9868 19892 9920
rect 19944 9908 19950 9920
rect 20714 9908 20720 9920
rect 19944 9880 20720 9908
rect 19944 9868 19950 9880
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 20824 9908 20852 9948
rect 21358 9936 21364 9988
rect 21416 9936 21422 9988
rect 21542 9908 21548 9920
rect 20824 9880 21548 9908
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 22204 9908 22232 10084
rect 23198 10072 23204 10124
rect 23256 10112 23262 10124
rect 23569 10115 23627 10121
rect 23569 10112 23581 10115
rect 23256 10084 23581 10112
rect 23256 10072 23262 10084
rect 23569 10081 23581 10084
rect 23615 10081 23627 10115
rect 23569 10075 23627 10081
rect 23661 10115 23719 10121
rect 23661 10081 23673 10115
rect 23707 10112 23719 10115
rect 24394 10112 24400 10124
rect 23707 10084 24400 10112
rect 23707 10081 23719 10084
rect 23661 10075 23719 10081
rect 24394 10072 24400 10084
rect 24452 10072 24458 10124
rect 24486 10072 24492 10124
rect 24544 10112 24550 10124
rect 24688 10112 24716 10152
rect 24544 10084 24716 10112
rect 24872 10112 24900 10152
rect 25590 10140 25596 10192
rect 25648 10180 25654 10192
rect 25685 10183 25743 10189
rect 25685 10180 25697 10183
rect 25648 10152 25697 10180
rect 25648 10140 25654 10152
rect 25685 10149 25697 10152
rect 25731 10180 25743 10183
rect 26510 10180 26516 10192
rect 25731 10152 26516 10180
rect 25731 10149 25743 10152
rect 25685 10143 25743 10149
rect 26510 10140 26516 10152
rect 26568 10140 26574 10192
rect 27080 10180 27108 10220
rect 30377 10217 30389 10220
rect 30423 10217 30435 10251
rect 30377 10211 30435 10217
rect 31662 10208 31668 10260
rect 31720 10208 31726 10260
rect 32398 10208 32404 10260
rect 32456 10248 32462 10260
rect 32674 10248 32680 10260
rect 32456 10220 32680 10248
rect 32456 10208 32462 10220
rect 32674 10208 32680 10220
rect 32732 10208 32738 10260
rect 32950 10208 32956 10260
rect 33008 10208 33014 10260
rect 33060 10220 36492 10248
rect 26712 10152 27108 10180
rect 26712 10112 26740 10152
rect 27154 10140 27160 10192
rect 27212 10180 27218 10192
rect 27614 10180 27620 10192
rect 27212 10152 27620 10180
rect 27212 10140 27218 10152
rect 27614 10140 27620 10152
rect 27672 10140 27678 10192
rect 27724 10152 29224 10180
rect 24872 10084 26740 10112
rect 24544 10072 24550 10084
rect 26786 10072 26792 10124
rect 26844 10112 26850 10124
rect 27724 10112 27752 10152
rect 26844 10084 27752 10112
rect 29196 10112 29224 10152
rect 29730 10140 29736 10192
rect 29788 10180 29794 10192
rect 31941 10183 31999 10189
rect 29788 10152 31708 10180
rect 29788 10140 29794 10152
rect 29196 10084 30972 10112
rect 26844 10072 26850 10084
rect 24785 10057 24843 10063
rect 22646 10004 22652 10056
rect 22704 10004 22710 10056
rect 23477 10047 23535 10053
rect 23477 10013 23489 10047
rect 23523 10044 23535 10047
rect 23750 10044 23756 10056
rect 23523 10016 23756 10044
rect 23523 10013 23535 10016
rect 23477 10007 23535 10013
rect 23750 10004 23756 10016
rect 23808 10004 23814 10056
rect 24673 10047 24731 10053
rect 24673 10013 24685 10047
rect 24719 10013 24731 10047
rect 24785 10023 24797 10057
rect 24831 10054 24843 10057
rect 24831 10026 24992 10054
rect 24831 10023 24843 10026
rect 24785 10017 24843 10023
rect 24673 10007 24731 10013
rect 24688 9976 24716 10007
rect 24762 9976 24768 9988
rect 24688 9948 24768 9976
rect 24762 9936 24768 9948
rect 24820 9936 24826 9988
rect 24964 9976 24992 10026
rect 25038 10004 25044 10056
rect 25096 10044 25102 10056
rect 26421 10047 26479 10053
rect 25096 10016 26372 10044
rect 25096 10004 25102 10016
rect 24964 9948 25084 9976
rect 25056 9920 25084 9948
rect 25682 9936 25688 9988
rect 25740 9936 25746 9988
rect 26142 9936 26148 9988
rect 26200 9936 26206 9988
rect 26344 9976 26372 10016
rect 26421 10013 26433 10047
rect 26467 10044 26479 10047
rect 26896 10044 27016 10046
rect 27614 10044 27620 10056
rect 26467 10018 27620 10044
rect 26467 10016 26924 10018
rect 26988 10016 27620 10018
rect 26467 10013 26479 10016
rect 26421 10007 26479 10013
rect 27614 10004 27620 10016
rect 27672 10004 27678 10056
rect 28350 10004 28356 10056
rect 28408 10044 28414 10056
rect 28537 10047 28595 10053
rect 28537 10044 28549 10047
rect 28408 10016 28549 10044
rect 28408 10004 28414 10016
rect 28537 10013 28549 10016
rect 28583 10013 28595 10047
rect 28537 10007 28595 10013
rect 28630 10047 28688 10053
rect 28630 10013 28642 10047
rect 28676 10013 28688 10047
rect 28630 10007 28688 10013
rect 26344 9948 26464 9976
rect 23109 9911 23167 9917
rect 23109 9908 23121 9911
rect 22204 9880 23121 9908
rect 23109 9877 23121 9880
rect 23155 9877 23167 9911
rect 23109 9871 23167 9877
rect 23750 9868 23756 9920
rect 23808 9908 23814 9920
rect 24949 9911 25007 9917
rect 24949 9908 24961 9911
rect 23808 9880 24961 9908
rect 23808 9868 23814 9880
rect 24949 9877 24961 9880
rect 24995 9877 25007 9911
rect 24949 9871 25007 9877
rect 25038 9868 25044 9920
rect 25096 9908 25102 9920
rect 25866 9908 25872 9920
rect 25096 9880 25872 9908
rect 25096 9868 25102 9880
rect 25866 9868 25872 9880
rect 25924 9868 25930 9920
rect 26234 9868 26240 9920
rect 26292 9868 26298 9920
rect 26436 9908 26464 9948
rect 27154 9936 27160 9988
rect 27212 9976 27218 9988
rect 27249 9979 27307 9985
rect 27249 9976 27261 9979
rect 27212 9948 27261 9976
rect 27212 9936 27218 9948
rect 27249 9945 27261 9948
rect 27295 9945 27307 9979
rect 27249 9939 27307 9945
rect 27430 9936 27436 9988
rect 27488 9936 27494 9988
rect 27522 9936 27528 9988
rect 27580 9936 27586 9988
rect 28258 9936 28264 9988
rect 28316 9976 28322 9988
rect 28645 9976 28673 10007
rect 28902 10006 28908 10058
rect 28960 10006 28966 10058
rect 29021 10047 29079 10053
rect 29021 10044 29033 10047
rect 29017 10013 29033 10044
rect 29067 10038 29079 10047
rect 29196 10038 29224 10084
rect 29067 10013 29224 10038
rect 29017 10010 29224 10013
rect 29733 10047 29791 10053
rect 29733 10013 29745 10047
rect 29779 10044 29791 10047
rect 30006 10044 30012 10056
rect 29779 10016 30012 10044
rect 29779 10013 29791 10016
rect 29021 10007 29079 10010
rect 29733 10007 29791 10013
rect 30006 10004 30012 10016
rect 30064 10004 30070 10056
rect 30742 10004 30748 10056
rect 30800 10004 30806 10056
rect 28813 9979 28871 9985
rect 28813 9976 28825 9979
rect 28316 9948 28673 9976
rect 28736 9948 28825 9976
rect 28316 9936 28322 9948
rect 27338 9908 27344 9920
rect 26436 9880 27344 9908
rect 27338 9868 27344 9880
rect 27396 9868 27402 9920
rect 28074 9868 28080 9920
rect 28132 9908 28138 9920
rect 28736 9908 28764 9948
rect 28813 9945 28825 9948
rect 28859 9945 28871 9979
rect 30944 9976 30972 10084
rect 31018 10072 31024 10124
rect 31076 10072 31082 10124
rect 31680 10121 31708 10152
rect 31941 10149 31953 10183
rect 31987 10180 31999 10183
rect 33060 10180 33088 10220
rect 36464 10180 36492 10220
rect 36538 10208 36544 10260
rect 36596 10248 36602 10260
rect 38565 10251 38623 10257
rect 38565 10248 38577 10251
rect 36596 10220 38577 10248
rect 36596 10208 36602 10220
rect 38565 10217 38577 10220
rect 38611 10217 38623 10251
rect 38565 10211 38623 10217
rect 36998 10180 37004 10192
rect 31987 10152 33088 10180
rect 33520 10152 33728 10180
rect 36464 10152 37004 10180
rect 31987 10149 31999 10152
rect 31941 10143 31999 10149
rect 31665 10115 31723 10121
rect 31665 10081 31677 10115
rect 31711 10081 31723 10115
rect 31665 10075 31723 10081
rect 32030 10072 32036 10124
rect 32088 10112 32094 10124
rect 33520 10112 33548 10152
rect 32088 10084 33548 10112
rect 32088 10072 32094 10084
rect 31573 10047 31631 10053
rect 31573 10013 31585 10047
rect 31619 10044 31631 10047
rect 31938 10044 31944 10056
rect 31619 10016 31944 10044
rect 31619 10013 31631 10016
rect 31573 10007 31631 10013
rect 31938 10004 31944 10016
rect 31996 10004 32002 10056
rect 32398 10004 32404 10056
rect 32456 10004 32462 10056
rect 32766 10044 32772 10056
rect 32508 10016 32772 10044
rect 32508 9976 32536 10016
rect 32766 10004 32772 10016
rect 32824 10004 32830 10056
rect 33410 10004 33416 10056
rect 33468 10004 33474 10056
rect 33700 10044 33728 10152
rect 36998 10140 37004 10152
rect 37056 10140 37062 10192
rect 34054 10072 34060 10124
rect 34112 10112 34118 10124
rect 34606 10112 34612 10124
rect 34112 10084 34612 10112
rect 34112 10072 34118 10084
rect 34606 10072 34612 10084
rect 34664 10112 34670 10124
rect 34885 10115 34943 10121
rect 34885 10112 34897 10115
rect 34664 10084 34897 10112
rect 34664 10072 34670 10084
rect 34885 10081 34897 10084
rect 34931 10081 34943 10115
rect 34885 10075 34943 10081
rect 33781 10047 33839 10053
rect 33781 10044 33793 10047
rect 33700 10016 33793 10044
rect 33781 10013 33793 10016
rect 33827 10013 33839 10047
rect 33962 10022 33968 10056
rect 33781 10007 33839 10013
rect 33904 10004 33968 10022
rect 34020 10004 34026 10056
rect 37369 10047 37427 10053
rect 37369 10013 37381 10047
rect 37415 10044 37427 10047
rect 37458 10044 37464 10056
rect 37415 10016 37464 10044
rect 37415 10013 37427 10016
rect 37369 10007 37427 10013
rect 37458 10004 37464 10016
rect 37516 10004 37522 10056
rect 38381 10047 38439 10053
rect 38381 10013 38393 10047
rect 38427 10044 38439 10047
rect 39390 10044 39396 10056
rect 38427 10016 39396 10044
rect 38427 10013 38439 10016
rect 38381 10007 38439 10013
rect 39390 10004 39396 10016
rect 39448 10004 39454 10056
rect 33904 9994 34008 10004
rect 30944 9948 32536 9976
rect 32585 9979 32643 9985
rect 28813 9939 28871 9945
rect 32585 9945 32597 9979
rect 32631 9945 32643 9979
rect 32585 9939 32643 9945
rect 32677 9979 32735 9985
rect 32677 9945 32689 9979
rect 32723 9976 32735 9979
rect 32858 9976 32864 9988
rect 32723 9948 32864 9976
rect 32723 9945 32735 9948
rect 32677 9939 32735 9945
rect 28132 9880 28764 9908
rect 29181 9911 29239 9917
rect 28132 9868 28138 9880
rect 29181 9877 29193 9911
rect 29227 9908 29239 9911
rect 29730 9908 29736 9920
rect 29227 9880 29736 9908
rect 29227 9877 29239 9880
rect 29181 9871 29239 9877
rect 29730 9868 29736 9880
rect 29788 9868 29794 9920
rect 29822 9868 29828 9920
rect 29880 9868 29886 9920
rect 30006 9868 30012 9920
rect 30064 9908 30070 9920
rect 30190 9908 30196 9920
rect 30064 9880 30196 9908
rect 30064 9868 30070 9880
rect 30190 9868 30196 9880
rect 30248 9868 30254 9920
rect 30837 9911 30895 9917
rect 30837 9877 30849 9911
rect 30883 9908 30895 9911
rect 31386 9908 31392 9920
rect 30883 9880 31392 9908
rect 30883 9877 30895 9880
rect 30837 9871 30895 9877
rect 31386 9868 31392 9880
rect 31444 9868 31450 9920
rect 31846 9868 31852 9920
rect 31904 9908 31910 9920
rect 32600 9908 32628 9939
rect 32858 9936 32864 9948
rect 32916 9936 32922 9988
rect 33597 9979 33655 9985
rect 33597 9945 33609 9979
rect 33643 9945 33655 9979
rect 33597 9939 33655 9945
rect 33689 9979 33747 9985
rect 33689 9945 33701 9979
rect 33735 9945 33747 9979
rect 33689 9939 33747 9945
rect 33612 9908 33640 9939
rect 31904 9880 33640 9908
rect 33704 9908 33732 9939
rect 33904 9908 33932 9994
rect 35158 9936 35164 9988
rect 35216 9936 35222 9988
rect 36446 9976 36452 9988
rect 36386 9948 36452 9976
rect 36446 9936 36452 9948
rect 36504 9936 36510 9988
rect 36909 9979 36967 9985
rect 36909 9945 36921 9979
rect 36955 9945 36967 9979
rect 36909 9939 36967 9945
rect 33704 9880 33932 9908
rect 31904 9868 31910 9880
rect 33962 9868 33968 9920
rect 34020 9868 34026 9920
rect 35342 9868 35348 9920
rect 35400 9908 35406 9920
rect 36924 9908 36952 9939
rect 35400 9880 36952 9908
rect 37461 9911 37519 9917
rect 35400 9868 35406 9880
rect 37461 9877 37473 9911
rect 37507 9908 37519 9911
rect 37550 9908 37556 9920
rect 37507 9880 37556 9908
rect 37507 9877 37519 9880
rect 37461 9871 37519 9877
rect 37550 9868 37556 9880
rect 37608 9868 37614 9920
rect 1104 9818 39352 9840
rect 1104 9766 10472 9818
rect 10524 9766 10536 9818
rect 10588 9766 10600 9818
rect 10652 9766 10664 9818
rect 10716 9766 10728 9818
rect 10780 9766 19994 9818
rect 20046 9766 20058 9818
rect 20110 9766 20122 9818
rect 20174 9766 20186 9818
rect 20238 9766 20250 9818
rect 20302 9766 29516 9818
rect 29568 9766 29580 9818
rect 29632 9766 29644 9818
rect 29696 9766 29708 9818
rect 29760 9766 29772 9818
rect 29824 9766 39038 9818
rect 39090 9766 39102 9818
rect 39154 9766 39166 9818
rect 39218 9766 39230 9818
rect 39282 9766 39294 9818
rect 39346 9766 39352 9818
rect 1104 9744 39352 9766
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 13633 9707 13691 9713
rect 13633 9704 13645 9707
rect 7156 9676 13645 9704
rect 7156 9664 7162 9676
rect 13633 9673 13645 9676
rect 13679 9673 13691 9707
rect 13633 9667 13691 9673
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 16114 9704 16120 9716
rect 13872 9676 16120 9704
rect 13872 9664 13878 9676
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 16482 9664 16488 9716
rect 16540 9704 16546 9716
rect 16850 9704 16856 9716
rect 16540 9676 16856 9704
rect 16540 9664 16546 9676
rect 16850 9664 16856 9676
rect 16908 9704 16914 9716
rect 17954 9704 17960 9716
rect 16908 9676 17960 9704
rect 16908 9664 16914 9676
rect 4893 9639 4951 9645
rect 4893 9636 4905 9639
rect 3910 9608 4905 9636
rect 4893 9605 4905 9608
rect 4939 9605 4951 9639
rect 5534 9636 5540 9648
rect 4893 9599 4951 9605
rect 5368 9608 5540 9636
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 1452 9540 1593 9568
rect 1452 9528 1458 9540
rect 1581 9537 1593 9540
rect 1627 9537 1639 9571
rect 1581 9531 1639 9537
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5368 9568 5396 9608
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 5629 9639 5687 9645
rect 5629 9605 5641 9639
rect 5675 9636 5687 9639
rect 6362 9636 6368 9648
rect 5675 9608 6368 9636
rect 5675 9605 5687 9608
rect 5629 9599 5687 9605
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 8754 9636 8760 9648
rect 8602 9608 8760 9636
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 9732 9608 10074 9636
rect 9732 9596 9738 9608
rect 11146 9596 11152 9648
rect 11204 9636 11210 9648
rect 11204 9608 12664 9636
rect 11204 9596 11210 9608
rect 4847 9540 5396 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 5442 9528 5448 9580
rect 5500 9528 5506 9580
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9537 5779 9571
rect 5721 9531 5779 9537
rect 2406 9460 2412 9512
rect 2464 9460 2470 9512
rect 2685 9503 2743 9509
rect 2685 9469 2697 9503
rect 2731 9500 2743 9503
rect 4154 9500 4160 9512
rect 2731 9472 4160 9500
rect 2731 9469 2743 9472
rect 2685 9463 2743 9469
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 5736 9500 5764 9531
rect 5810 9528 5816 9580
rect 5868 9528 5874 9580
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9568 11851 9571
rect 11974 9568 11980 9580
rect 11839 9540 11980 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12526 9528 12532 9580
rect 12584 9528 12590 9580
rect 12636 9568 12664 9608
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 14093 9639 14151 9645
rect 14093 9636 14105 9639
rect 12768 9608 14105 9636
rect 12768 9596 12774 9608
rect 14093 9605 14105 9608
rect 14139 9605 14151 9639
rect 14093 9599 14151 9605
rect 15197 9639 15255 9645
rect 15197 9605 15209 9639
rect 15243 9636 15255 9639
rect 15243 9608 16068 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 13906 9568 13912 9580
rect 12636 9540 13912 9568
rect 13906 9528 13912 9540
rect 13964 9568 13970 9580
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 13964 9540 14013 9568
rect 13964 9528 13970 9540
rect 14001 9537 14013 9540
rect 14047 9537 14059 9571
rect 14458 9568 14464 9580
rect 14001 9531 14059 9537
rect 14292 9540 14464 9568
rect 4304 9472 5764 9500
rect 4304 9460 4310 9472
rect 6270 9460 6276 9512
rect 6328 9500 6334 9512
rect 6822 9500 6828 9512
rect 6328 9472 6828 9500
rect 6328 9460 6334 9472
rect 6822 9460 6828 9472
rect 6880 9500 6886 9512
rect 7101 9503 7159 9509
rect 7101 9500 7113 9503
rect 6880 9472 7113 9500
rect 6880 9460 6886 9472
rect 7101 9469 7113 9472
rect 7147 9469 7159 9503
rect 7101 9463 7159 9469
rect 7374 9460 7380 9512
rect 7432 9460 7438 9512
rect 8110 9460 8116 9512
rect 8168 9500 8174 9512
rect 9306 9500 9312 9512
rect 8168 9472 9312 9500
rect 8168 9460 8174 9472
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 9582 9460 9588 9512
rect 9640 9460 9646 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 11606 9500 11612 9512
rect 9732 9472 11612 9500
rect 9732 9460 9738 9472
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 11940 9472 13093 9500
rect 11940 9460 11946 9472
rect 13081 9469 13093 9472
rect 13127 9500 13139 9503
rect 13170 9500 13176 9512
rect 13127 9472 13176 9500
rect 13127 9469 13139 9472
rect 13081 9463 13139 9469
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 14292 9509 14320 9540
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 14700 9540 15240 9568
rect 14700 9528 14706 9540
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9469 14335 9503
rect 15102 9500 15108 9512
rect 14277 9463 14335 9469
rect 14384 9472 15108 9500
rect 4080 9404 7236 9432
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 4080 9364 4108 9404
rect 7208 9376 7236 9404
rect 8478 9392 8484 9444
rect 8536 9432 8542 9444
rect 8754 9432 8760 9444
rect 8536 9404 8760 9432
rect 8536 9392 8542 9404
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 10594 9392 10600 9444
rect 10652 9432 10658 9444
rect 11057 9435 11115 9441
rect 11057 9432 11069 9435
rect 10652 9404 11069 9432
rect 10652 9392 10658 9404
rect 11057 9401 11069 9404
rect 11103 9432 11115 9435
rect 12066 9432 12072 9444
rect 11103 9404 12072 9432
rect 11103 9401 11115 9404
rect 11057 9395 11115 9401
rect 12066 9392 12072 9404
rect 12124 9392 12130 9444
rect 12710 9392 12716 9444
rect 12768 9432 12774 9444
rect 14384 9432 14412 9472
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 15212 9500 15240 9540
rect 15286 9528 15292 9580
rect 15344 9528 15350 9580
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 15212 9472 15393 9500
rect 15381 9469 15393 9472
rect 15427 9469 15439 9503
rect 16040 9500 16068 9608
rect 16206 9596 16212 9648
rect 16264 9596 16270 9648
rect 17034 9596 17040 9648
rect 17092 9636 17098 9648
rect 17589 9639 17647 9645
rect 17589 9636 17601 9639
rect 17092 9608 17601 9636
rect 17092 9596 17098 9608
rect 17589 9605 17601 9608
rect 17635 9605 17647 9639
rect 17589 9599 17647 9605
rect 17770 9596 17776 9648
rect 17828 9596 17834 9648
rect 17880 9645 17908 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 19886 9664 19892 9716
rect 19944 9704 19950 9716
rect 20806 9704 20812 9716
rect 19944 9676 20812 9704
rect 19944 9664 19950 9676
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 22646 9704 22652 9716
rect 21652 9676 22652 9704
rect 17865 9639 17923 9645
rect 17865 9605 17877 9639
rect 17911 9605 17923 9639
rect 17865 9599 17923 9605
rect 20346 9596 20352 9648
rect 20404 9636 20410 9648
rect 21177 9639 21235 9645
rect 21177 9636 21189 9639
rect 20404 9608 21189 9636
rect 20404 9596 20410 9608
rect 21177 9605 21189 9608
rect 21223 9605 21235 9639
rect 21177 9599 21235 9605
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 16298 9568 16304 9580
rect 16163 9540 16304 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 16298 9528 16304 9540
rect 16356 9568 16362 9580
rect 16482 9568 16488 9580
rect 16356 9540 16488 9568
rect 16356 9528 16362 9540
rect 16482 9528 16488 9540
rect 16540 9528 16546 9580
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 18693 9571 18751 9577
rect 18693 9568 18705 9571
rect 16816 9540 18705 9568
rect 16816 9528 16822 9540
rect 17880 9512 17908 9540
rect 18693 9537 18705 9540
rect 18739 9537 18751 9571
rect 20438 9568 20444 9580
rect 20102 9540 20444 9568
rect 18693 9531 18751 9537
rect 20438 9528 20444 9540
rect 20496 9528 20502 9580
rect 20901 9571 20959 9577
rect 20901 9537 20913 9571
rect 20947 9568 20959 9571
rect 20990 9568 20996 9580
rect 20947 9540 20996 9568
rect 20947 9537 20959 9540
rect 20901 9531 20959 9537
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 21085 9571 21143 9577
rect 21085 9537 21097 9571
rect 21131 9537 21143 9571
rect 21085 9531 21143 9537
rect 17586 9500 17592 9512
rect 16040 9472 17592 9500
rect 15381 9463 15439 9469
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 17862 9460 17868 9512
rect 17920 9460 17926 9512
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 17972 9472 18981 9500
rect 12768 9404 14412 9432
rect 14829 9435 14887 9441
rect 12768 9392 12774 9404
rect 14829 9401 14841 9435
rect 14875 9401 14887 9435
rect 14829 9395 14887 9401
rect 1811 9336 4108 9364
rect 4157 9367 4215 9373
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4522 9364 4528 9376
rect 4203 9336 4528 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4522 9324 4528 9336
rect 4580 9364 4586 9376
rect 5534 9364 5540 9376
rect 4580 9336 5540 9364
rect 4580 9324 4586 9336
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5997 9367 6055 9373
rect 5997 9333 6009 9367
rect 6043 9364 6055 9367
rect 6086 9364 6092 9376
rect 6043 9336 6092 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 7190 9324 7196 9376
rect 7248 9324 7254 9376
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 7616 9336 8861 9364
rect 7616 9324 7622 9336
rect 8849 9333 8861 9336
rect 8895 9333 8907 9367
rect 8849 9327 8907 9333
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 11698 9364 11704 9376
rect 8996 9336 11704 9364
rect 8996 9324 9002 9336
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 11882 9324 11888 9376
rect 11940 9324 11946 9376
rect 14844 9364 14872 9395
rect 15470 9392 15476 9444
rect 15528 9432 15534 9444
rect 16206 9432 16212 9444
rect 15528 9404 16212 9432
rect 15528 9392 15534 9404
rect 16206 9392 16212 9404
rect 16264 9392 16270 9444
rect 17972 9432 18000 9472
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 19702 9460 19708 9512
rect 19760 9500 19766 9512
rect 21100 9500 21128 9531
rect 21266 9528 21272 9580
rect 21324 9568 21330 9580
rect 21652 9568 21680 9676
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 26510 9704 26516 9716
rect 26482 9664 26516 9704
rect 26568 9704 26574 9716
rect 26568 9676 26740 9704
rect 26568 9664 26574 9676
rect 22097 9639 22155 9645
rect 22097 9605 22109 9639
rect 22143 9636 22155 9639
rect 22554 9636 22560 9648
rect 22143 9608 22560 9636
rect 22143 9605 22155 9608
rect 22097 9599 22155 9605
rect 22554 9596 22560 9608
rect 22612 9596 22618 9648
rect 23934 9636 23940 9648
rect 23584 9608 23940 9636
rect 21324 9540 21680 9568
rect 22244 9571 22302 9577
rect 21324 9528 21330 9540
rect 22244 9537 22256 9571
rect 22290 9568 22302 9571
rect 23584 9568 23612 9608
rect 23934 9596 23940 9608
rect 23992 9596 23998 9648
rect 24026 9596 24032 9648
rect 24084 9596 24090 9648
rect 25314 9596 25320 9648
rect 25372 9636 25378 9648
rect 25372 9608 26280 9636
rect 25372 9596 25378 9608
rect 22290 9540 23612 9568
rect 22290 9537 22302 9540
rect 22244 9531 22302 9537
rect 23658 9528 23664 9580
rect 23716 9568 23722 9580
rect 23753 9571 23811 9577
rect 23753 9568 23765 9571
rect 23716 9540 23765 9568
rect 23716 9528 23722 9540
rect 23753 9537 23765 9540
rect 23799 9537 23811 9571
rect 23753 9531 23811 9537
rect 25130 9528 25136 9580
rect 25188 9528 25194 9580
rect 25682 9528 25688 9580
rect 25740 9568 25746 9580
rect 26252 9577 26280 9608
rect 26482 9602 26510 9664
rect 26436 9577 26510 9602
rect 26712 9580 26740 9676
rect 27586 9676 29045 9704
rect 26786 9596 26792 9648
rect 26844 9636 26850 9648
rect 27586 9636 27614 9676
rect 26844 9608 27614 9636
rect 26844 9596 26850 9608
rect 27890 9596 27896 9648
rect 27948 9596 27954 9648
rect 27982 9596 27988 9648
rect 28040 9596 28046 9648
rect 28813 9639 28871 9645
rect 28813 9636 28825 9639
rect 28097 9608 28825 9636
rect 26053 9571 26111 9577
rect 26053 9568 26065 9571
rect 25740 9540 26065 9568
rect 25740 9528 25746 9540
rect 26053 9537 26065 9540
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 26237 9571 26295 9577
rect 26237 9537 26249 9571
rect 26283 9537 26295 9571
rect 26237 9531 26295 9537
rect 26329 9571 26387 9577
rect 26329 9537 26341 9571
rect 26375 9537 26387 9571
rect 26329 9531 26387 9537
rect 26421 9574 26510 9577
rect 26421 9571 26479 9574
rect 26421 9537 26433 9571
rect 26467 9537 26479 9571
rect 26421 9531 26479 9537
rect 22465 9503 22523 9509
rect 19760 9472 22232 9500
rect 19760 9460 19766 9472
rect 16684 9404 18000 9432
rect 21453 9435 21511 9441
rect 16684 9364 16712 9404
rect 21453 9401 21465 9435
rect 21499 9432 21511 9435
rect 22204 9432 22232 9472
rect 22465 9469 22477 9503
rect 22511 9500 22523 9503
rect 22511 9472 22692 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 22664 9432 22692 9472
rect 22738 9460 22744 9512
rect 22796 9460 22802 9512
rect 23750 9432 23756 9444
rect 21499 9404 22094 9432
rect 22204 9404 22495 9432
rect 22664 9404 23756 9432
rect 21499 9401 21511 9404
rect 21453 9395 21511 9401
rect 14844 9336 16712 9364
rect 17310 9324 17316 9376
rect 17368 9324 17374 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 20441 9367 20499 9373
rect 20441 9364 20453 9367
rect 18288 9336 20453 9364
rect 18288 9324 18294 9336
rect 20441 9333 20453 9336
rect 20487 9333 20499 9367
rect 22066 9364 22094 9404
rect 22373 9367 22431 9373
rect 22373 9364 22385 9367
rect 22066 9336 22385 9364
rect 20441 9327 20499 9333
rect 22373 9333 22385 9336
rect 22419 9333 22431 9367
rect 22467 9364 22495 9404
rect 23750 9392 23756 9404
rect 23808 9392 23814 9444
rect 26142 9392 26148 9444
rect 26200 9432 26206 9444
rect 26344 9432 26372 9531
rect 26694 9528 26700 9580
rect 26752 9568 26758 9580
rect 26752 9540 27844 9568
rect 26752 9528 26758 9540
rect 27522 9500 27528 9512
rect 26528 9472 27528 9500
rect 26528 9444 26556 9472
rect 27522 9460 27528 9472
rect 27580 9500 27586 9512
rect 27816 9500 27844 9540
rect 27890 9500 27896 9512
rect 27580 9472 27667 9500
rect 27816 9472 27896 9500
rect 27580 9460 27586 9472
rect 26200 9404 26372 9432
rect 26200 9392 26206 9404
rect 26510 9392 26516 9444
rect 26568 9392 26574 9444
rect 26605 9435 26663 9441
rect 26605 9401 26617 9435
rect 26651 9432 26663 9435
rect 27154 9432 27160 9444
rect 26651 9404 27160 9432
rect 26651 9401 26663 9404
rect 26605 9395 26663 9401
rect 27154 9392 27160 9404
rect 27212 9392 27218 9444
rect 25314 9364 25320 9376
rect 22467 9336 25320 9364
rect 22373 9327 22431 9333
rect 25314 9324 25320 9336
rect 25372 9324 25378 9376
rect 25498 9324 25504 9376
rect 25556 9324 25562 9376
rect 25590 9324 25596 9376
rect 25648 9364 25654 9376
rect 26786 9364 26792 9376
rect 25648 9336 26792 9364
rect 25648 9324 25654 9336
rect 26786 9324 26792 9336
rect 26844 9324 26850 9376
rect 27430 9324 27436 9376
rect 27488 9364 27494 9376
rect 27525 9367 27583 9373
rect 27525 9364 27537 9367
rect 27488 9336 27537 9364
rect 27488 9324 27494 9336
rect 27525 9333 27537 9336
rect 27571 9333 27583 9367
rect 27639 9364 27667 9472
rect 27890 9460 27896 9472
rect 27948 9460 27954 9512
rect 27706 9392 27712 9444
rect 27764 9432 27770 9444
rect 28097 9432 28125 9608
rect 28813 9605 28825 9608
rect 28859 9605 28871 9639
rect 29017 9636 29045 9676
rect 29086 9664 29092 9716
rect 29144 9704 29150 9716
rect 29273 9707 29331 9713
rect 29273 9704 29285 9707
rect 29144 9676 29285 9704
rect 29144 9664 29150 9676
rect 29273 9673 29285 9676
rect 29319 9673 29331 9707
rect 29273 9667 29331 9673
rect 29365 9707 29423 9713
rect 29365 9673 29377 9707
rect 29411 9704 29423 9707
rect 29454 9704 29460 9716
rect 29411 9676 29460 9704
rect 29411 9673 29423 9676
rect 29365 9667 29423 9673
rect 29454 9664 29460 9676
rect 29512 9664 29518 9716
rect 29546 9664 29552 9716
rect 29604 9704 29610 9716
rect 30282 9704 30288 9716
rect 29604 9676 30288 9704
rect 29604 9664 29610 9676
rect 30282 9664 30288 9676
rect 30340 9664 30346 9716
rect 31018 9704 31024 9716
rect 30668 9676 31024 9704
rect 29178 9636 29184 9648
rect 29017 9608 29184 9636
rect 28813 9599 28871 9605
rect 29178 9596 29184 9608
rect 29236 9596 29242 9648
rect 30668 9636 30696 9676
rect 31018 9664 31024 9676
rect 31076 9704 31082 9716
rect 31662 9704 31668 9716
rect 31076 9676 31668 9704
rect 31076 9664 31082 9676
rect 31662 9664 31668 9676
rect 31720 9704 31726 9716
rect 33042 9704 33048 9716
rect 31720 9676 33048 9704
rect 31720 9664 31726 9676
rect 33042 9664 33048 9676
rect 33100 9664 33106 9716
rect 33428 9676 34836 9704
rect 33428 9636 33456 9676
rect 30024 9608 30696 9636
rect 31772 9608 33456 9636
rect 33505 9639 33563 9645
rect 28276 9568 28488 9574
rect 30024 9568 30052 9608
rect 28276 9546 30052 9568
rect 28169 9503 28227 9509
rect 28169 9469 28181 9503
rect 28215 9500 28227 9503
rect 28276 9500 28304 9546
rect 28460 9540 30052 9546
rect 28215 9472 28304 9500
rect 28215 9469 28227 9472
rect 28169 9463 28227 9469
rect 28350 9460 28356 9512
rect 28408 9500 28414 9512
rect 29549 9503 29607 9509
rect 29549 9500 29561 9503
rect 28408 9472 29561 9500
rect 28408 9460 28414 9472
rect 29549 9469 29561 9472
rect 29595 9469 29607 9503
rect 29549 9463 29607 9469
rect 30006 9460 30012 9512
rect 30064 9460 30070 9512
rect 30285 9503 30343 9509
rect 30285 9469 30297 9503
rect 30331 9500 30343 9503
rect 31018 9500 31024 9512
rect 30331 9472 31024 9500
rect 30331 9469 30343 9472
rect 30285 9463 30343 9469
rect 31018 9460 31024 9472
rect 31076 9460 31082 9512
rect 28813 9435 28871 9441
rect 27764 9404 28125 9432
rect 28368 9404 28764 9432
rect 27764 9392 27770 9404
rect 28368 9364 28396 9404
rect 27639 9336 28396 9364
rect 28736 9364 28764 9404
rect 28813 9401 28825 9435
rect 28859 9432 28871 9435
rect 29178 9432 29184 9444
rect 28859 9404 29184 9432
rect 28859 9401 28871 9404
rect 28813 9395 28871 9401
rect 29178 9392 29184 9404
rect 29236 9392 29242 9444
rect 31404 9432 31432 9554
rect 31772 9509 31800 9608
rect 33505 9605 33517 9639
rect 33551 9636 33563 9639
rect 33778 9636 33784 9648
rect 33551 9608 33784 9636
rect 33551 9605 33563 9608
rect 33505 9599 33563 9605
rect 33778 9596 33784 9608
rect 33836 9596 33842 9648
rect 34514 9596 34520 9648
rect 34572 9596 34578 9648
rect 34808 9636 34836 9676
rect 34808 9608 36124 9636
rect 31938 9528 31944 9580
rect 31996 9568 32002 9580
rect 32309 9571 32367 9577
rect 32309 9568 32321 9571
rect 31996 9540 32321 9568
rect 31996 9528 32002 9540
rect 32309 9537 32321 9540
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 35618 9528 35624 9580
rect 35676 9528 35682 9580
rect 31757 9503 31815 9509
rect 31757 9469 31769 9503
rect 31803 9469 31815 9503
rect 31757 9463 31815 9469
rect 32582 9460 32588 9512
rect 32640 9460 32646 9512
rect 33226 9460 33232 9512
rect 33284 9460 33290 9512
rect 36096 9500 36124 9608
rect 36538 9596 36544 9648
rect 36596 9636 36602 9648
rect 36817 9639 36875 9645
rect 36817 9636 36829 9639
rect 36596 9608 36829 9636
rect 36596 9596 36602 9608
rect 36817 9605 36829 9608
rect 36863 9605 36875 9639
rect 36817 9599 36875 9605
rect 36173 9571 36231 9577
rect 36173 9537 36185 9571
rect 36219 9568 36231 9571
rect 36725 9571 36783 9577
rect 36725 9568 36737 9571
rect 36219 9540 36737 9568
rect 36219 9537 36231 9540
rect 36173 9531 36231 9537
rect 36725 9537 36737 9540
rect 36771 9568 36783 9571
rect 37458 9568 37464 9580
rect 36771 9540 37464 9568
rect 36771 9537 36783 9540
rect 36725 9531 36783 9537
rect 37458 9528 37464 9540
rect 37516 9528 37522 9580
rect 38102 9528 38108 9580
rect 38160 9528 38166 9580
rect 37918 9500 37924 9512
rect 33336 9472 34560 9500
rect 36096 9472 37924 9500
rect 33336 9432 33364 9472
rect 31404 9404 33364 9432
rect 34532 9432 34560 9472
rect 37918 9460 37924 9472
rect 37976 9460 37982 9512
rect 37553 9435 37611 9441
rect 37553 9432 37565 9435
rect 34532 9404 37565 9432
rect 37553 9401 37565 9404
rect 37599 9401 37611 9435
rect 37553 9395 37611 9401
rect 31478 9364 31484 9376
rect 28736 9336 31484 9364
rect 27525 9327 27583 9333
rect 31478 9324 31484 9336
rect 31536 9324 31542 9376
rect 33318 9324 33324 9376
rect 33376 9364 33382 9376
rect 34977 9367 35035 9373
rect 34977 9364 34989 9367
rect 33376 9336 34989 9364
rect 33376 9324 33382 9336
rect 34977 9333 34989 9336
rect 35023 9333 35035 9367
rect 34977 9327 35035 9333
rect 38194 9324 38200 9376
rect 38252 9324 38258 9376
rect 1104 9274 39192 9296
rect 1104 9222 5711 9274
rect 5763 9222 5775 9274
rect 5827 9222 5839 9274
rect 5891 9222 5903 9274
rect 5955 9222 5967 9274
rect 6019 9222 15233 9274
rect 15285 9222 15297 9274
rect 15349 9222 15361 9274
rect 15413 9222 15425 9274
rect 15477 9222 15489 9274
rect 15541 9222 24755 9274
rect 24807 9222 24819 9274
rect 24871 9222 24883 9274
rect 24935 9222 24947 9274
rect 24999 9222 25011 9274
rect 25063 9222 34277 9274
rect 34329 9222 34341 9274
rect 34393 9222 34405 9274
rect 34457 9222 34469 9274
rect 34521 9222 34533 9274
rect 34585 9222 39192 9274
rect 1104 9200 39192 9222
rect 2314 9120 2320 9172
rect 2372 9120 2378 9172
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 4062 9160 4068 9172
rect 3016 9132 4068 9160
rect 3016 9120 3022 9132
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4236 9163 4294 9169
rect 4236 9129 4248 9163
rect 4282 9160 4294 9163
rect 5994 9160 6000 9172
rect 4282 9132 6000 9160
rect 4282 9129 4294 9132
rect 4236 9123 4294 9129
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9160 6607 9163
rect 7374 9160 7380 9172
rect 6595 9132 7380 9160
rect 6595 9129 6607 9132
rect 6549 9123 6607 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8202 9160 8208 9172
rect 7800 9132 8208 9160
rect 7800 9120 7806 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8386 9120 8392 9172
rect 8444 9120 8450 9172
rect 9401 9163 9459 9169
rect 9401 9129 9413 9163
rect 9447 9160 9459 9163
rect 9582 9160 9588 9172
rect 9447 9132 9588 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 12805 9163 12863 9169
rect 12805 9160 12817 9163
rect 11992 9132 12817 9160
rect 2406 9052 2412 9104
rect 2464 9092 2470 9104
rect 2464 9064 4016 9092
rect 2464 9052 2470 9064
rect 2130 8984 2136 9036
rect 2188 9024 2194 9036
rect 2590 9024 2596 9036
rect 2188 8996 2596 9024
rect 2188 8984 2194 8996
rect 2590 8984 2596 8996
rect 2648 9024 2654 9036
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2648 8996 2881 9024
rect 2648 8984 2654 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 3694 9024 3700 9036
rect 3200 8996 3700 9024
rect 3200 8984 3206 8996
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 3988 9033 4016 9064
rect 6086 9052 6092 9104
rect 6144 9092 6150 9104
rect 8938 9092 8944 9104
rect 6144 9064 8944 9092
rect 6144 9052 6150 9064
rect 8938 9052 8944 9064
rect 8996 9052 9002 9104
rect 11992 9092 12020 9132
rect 12805 9129 12817 9132
rect 12851 9129 12863 9163
rect 12805 9123 12863 9129
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 15562 9160 15568 9172
rect 14792 9132 15568 9160
rect 14792 9120 14798 9132
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 22370 9160 22376 9172
rect 18616 9132 22376 9160
rect 11900 9064 12020 9092
rect 12345 9095 12403 9101
rect 3973 9027 4031 9033
rect 3973 8993 3985 9027
rect 4019 9024 4031 9027
rect 4246 9024 4252 9036
rect 4019 8996 4252 9024
rect 4019 8993 4031 8996
rect 3973 8987 4031 8993
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 4798 8984 4804 9036
rect 4856 9024 4862 9036
rect 7098 9024 7104 9036
rect 4856 8996 7104 9024
rect 4856 8984 4862 8996
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 9674 9024 9680 9036
rect 7760 8996 9680 9024
rect 14 8916 20 8968
rect 72 8956 78 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 72 8928 1593 8956
rect 72 8916 78 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 3786 8956 3792 8968
rect 2731 8928 3792 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 5684 8928 6929 8956
rect 5684 8916 5690 8928
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8956 7067 8959
rect 7558 8956 7564 8968
rect 7055 8928 7564 8956
rect 7055 8925 7067 8928
rect 7009 8919 7067 8925
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 7760 8965 7788 8996
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10318 9024 10324 9036
rect 10091 8996 10324 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 9024 10655 9027
rect 10962 9024 10968 9036
rect 10643 8996 10968 9024
rect 10643 8993 10655 8996
rect 10597 8987 10655 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11900 9024 11928 9064
rect 12345 9061 12357 9095
rect 12391 9092 12403 9095
rect 12526 9092 12532 9104
rect 12391 9064 12532 9092
rect 12391 9061 12403 9064
rect 12345 9055 12403 9061
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 13372 9064 13584 9092
rect 13372 9024 13400 9064
rect 11388 8996 11928 9024
rect 12268 8996 13400 9024
rect 11388 8984 11394 8996
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7834 8916 7840 8968
rect 7892 8916 7898 8968
rect 7926 8916 7932 8968
rect 7984 8956 7990 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 7984 8928 8125 8956
rect 7984 8916 7990 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 8202 8916 8208 8968
rect 8260 8965 8266 8968
rect 8260 8956 8268 8965
rect 9769 8959 9827 8965
rect 8260 8928 8305 8956
rect 8260 8919 8268 8928
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 10410 8956 10416 8968
rect 9815 8928 10416 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 8260 8916 8266 8919
rect 2777 8891 2835 8897
rect 2777 8857 2789 8891
rect 2823 8888 2835 8891
rect 2823 8860 2857 8888
rect 2823 8857 2835 8860
rect 2777 8851 2835 8857
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8820 1823 8823
rect 2792 8820 2820 8851
rect 4982 8848 4988 8900
rect 5040 8848 5046 8900
rect 6362 8848 6368 8900
rect 6420 8888 6426 8900
rect 6420 8860 7881 8888
rect 6420 8848 6426 8860
rect 5074 8820 5080 8832
rect 1811 8792 5080 8820
rect 1811 8789 1823 8792
rect 1765 8783 1823 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5721 8823 5779 8829
rect 5721 8789 5733 8823
rect 5767 8820 5779 8823
rect 6822 8820 6828 8832
rect 5767 8792 6828 8820
rect 5767 8789 5779 8792
rect 5721 8783 5779 8789
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7190 8780 7196 8832
rect 7248 8820 7254 8832
rect 7742 8820 7748 8832
rect 7248 8792 7748 8820
rect 7248 8780 7254 8792
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 7853 8820 7881 8860
rect 8018 8848 8024 8900
rect 8076 8848 8082 8900
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 9784 8888 9812 8919
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 9732 8860 9812 8888
rect 9861 8891 9919 8897
rect 9732 8848 9738 8860
rect 9861 8857 9873 8891
rect 9907 8888 9919 8891
rect 10594 8888 10600 8900
rect 9907 8860 10600 8888
rect 9907 8857 9919 8860
rect 9861 8851 9919 8857
rect 10594 8848 10600 8860
rect 10652 8848 10658 8900
rect 10873 8891 10931 8897
rect 10873 8857 10885 8891
rect 10919 8857 10931 8891
rect 10873 8851 10931 8857
rect 10778 8820 10784 8832
rect 7853 8792 10784 8820
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 10888 8820 10916 8851
rect 11882 8848 11888 8900
rect 11940 8848 11946 8900
rect 12268 8820 12296 8996
rect 13446 8984 13452 9036
rect 13504 8984 13510 9036
rect 13556 9024 13584 9064
rect 14458 9052 14464 9104
rect 14516 9092 14522 9104
rect 14826 9092 14832 9104
rect 14516 9064 14832 9092
rect 14516 9052 14522 9064
rect 14826 9052 14832 9064
rect 14884 9052 14890 9104
rect 15212 9064 15608 9092
rect 13906 9024 13912 9036
rect 13556 8996 13912 9024
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 14182 8984 14188 9036
rect 14240 9024 14246 9036
rect 14938 9027 14996 9033
rect 14240 8996 14688 9024
rect 14240 8984 14246 8996
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 14274 8956 14280 8968
rect 13219 8928 14280 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 14366 8916 14372 8968
rect 14424 8916 14430 8968
rect 12894 8848 12900 8900
rect 12952 8888 12958 8900
rect 14660 8897 14688 8996
rect 14938 8993 14950 9027
rect 14984 9024 14996 9027
rect 15102 9024 15108 9036
rect 14984 8996 15108 9024
rect 14984 8993 14996 8996
rect 14938 8987 14996 8993
rect 15102 8984 15108 8996
rect 15160 8984 15166 9036
rect 14826 8965 14832 8968
rect 14789 8959 14832 8965
rect 14789 8925 14801 8959
rect 14884 8956 14890 8968
rect 15212 8956 15240 9064
rect 15470 8984 15476 9036
rect 15528 8984 15534 9036
rect 15580 9024 15608 9064
rect 15838 9024 15844 9036
rect 15580 8996 15844 9024
rect 15838 8984 15844 8996
rect 15896 9024 15902 9036
rect 15896 8996 17264 9024
rect 15896 8984 15902 8996
rect 14884 8928 15240 8956
rect 14789 8919 14832 8925
rect 14826 8916 14832 8919
rect 14884 8916 14890 8928
rect 13265 8891 13323 8897
rect 13265 8888 13277 8891
rect 12952 8860 13277 8888
rect 12952 8848 12958 8860
rect 13265 8857 13277 8860
rect 13311 8857 13323 8891
rect 13265 8851 13323 8857
rect 14553 8891 14611 8897
rect 14553 8857 14565 8891
rect 14599 8857 14611 8891
rect 14553 8851 14611 8857
rect 14645 8891 14703 8897
rect 14645 8857 14657 8891
rect 14691 8857 14703 8891
rect 15378 8888 15384 8900
rect 14645 8851 14703 8857
rect 15212 8860 15384 8888
rect 10888 8792 12296 8820
rect 13630 8780 13636 8832
rect 13688 8820 13694 8832
rect 14568 8820 14596 8851
rect 13688 8792 14596 8820
rect 13688 8780 13694 8792
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 15212 8820 15240 8860
rect 15378 8848 15384 8860
rect 15436 8848 15442 8900
rect 15746 8848 15752 8900
rect 15804 8848 15810 8900
rect 15856 8860 16238 8888
rect 14792 8792 15240 8820
rect 14792 8780 14798 8792
rect 15286 8780 15292 8832
rect 15344 8820 15350 8832
rect 15856 8820 15884 8860
rect 15344 8792 15884 8820
rect 17236 8820 17264 8996
rect 17586 8916 17592 8968
rect 17644 8956 17650 8968
rect 18230 8956 18236 8968
rect 17644 8928 18236 8956
rect 17644 8916 17650 8928
rect 18230 8916 18236 8928
rect 18288 8956 18294 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 18288 8928 18337 8956
rect 18288 8916 18294 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8956 18567 8959
rect 18616 8956 18644 9132
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 25590 9160 25596 9172
rect 22848 9132 25596 9160
rect 22848 9101 22876 9132
rect 25590 9120 25596 9132
rect 25648 9120 25654 9172
rect 26234 9120 26240 9172
rect 26292 9160 26298 9172
rect 26329 9163 26387 9169
rect 26329 9160 26341 9163
rect 26292 9132 26341 9160
rect 26292 9120 26298 9132
rect 26329 9129 26341 9132
rect 26375 9129 26387 9163
rect 26329 9123 26387 9129
rect 26418 9120 26424 9172
rect 26476 9160 26482 9172
rect 26602 9160 26608 9172
rect 26476 9132 26608 9160
rect 26476 9120 26482 9132
rect 26602 9120 26608 9132
rect 26660 9120 26666 9172
rect 30742 9160 30748 9172
rect 27356 9132 30748 9160
rect 22833 9095 22891 9101
rect 19260 9064 20668 9092
rect 18555 8928 18644 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 18690 8916 18696 8968
rect 18748 8916 18754 8968
rect 19260 8956 19288 9064
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19392 8996 19565 9024
rect 19392 8984 19398 8996
rect 19537 8965 19565 8996
rect 20530 8984 20536 9036
rect 20588 8984 20594 9036
rect 20640 9024 20668 9064
rect 22833 9061 22845 9095
rect 22879 9061 22891 9095
rect 27356 9092 27384 9132
rect 30742 9120 30748 9132
rect 30800 9120 30806 9172
rect 31018 9120 31024 9172
rect 31076 9160 31082 9172
rect 34698 9160 34704 9172
rect 31076 9132 34704 9160
rect 31076 9120 31082 9132
rect 34698 9120 34704 9132
rect 34756 9120 34762 9172
rect 34885 9163 34943 9169
rect 34885 9129 34897 9163
rect 34931 9160 34943 9163
rect 35158 9160 35164 9172
rect 34931 9132 35164 9160
rect 34931 9129 34943 9132
rect 34885 9123 34943 9129
rect 35158 9120 35164 9132
rect 35216 9120 35222 9172
rect 36170 9120 36176 9172
rect 36228 9120 36234 9172
rect 38562 9120 38568 9172
rect 38620 9120 38626 9172
rect 22833 9055 22891 9061
rect 26436 9064 27384 9092
rect 28997 9095 29055 9101
rect 26436 9036 26464 9064
rect 28997 9061 29009 9095
rect 29043 9092 29055 9095
rect 29270 9092 29276 9104
rect 29043 9064 29276 9092
rect 29043 9061 29055 9064
rect 28997 9055 29055 9061
rect 29270 9052 29276 9064
rect 29328 9052 29334 9104
rect 30190 9052 30196 9104
rect 30248 9092 30254 9104
rect 30285 9095 30343 9101
rect 30285 9092 30297 9095
rect 30248 9064 30297 9092
rect 30248 9052 30254 9064
rect 30285 9061 30297 9064
rect 30331 9061 30343 9095
rect 30285 9055 30343 9061
rect 32582 9052 32588 9104
rect 32640 9092 32646 9104
rect 34606 9092 34612 9104
rect 32640 9064 34612 9092
rect 32640 9052 32646 9064
rect 34606 9052 34612 9064
rect 34664 9092 34670 9104
rect 35618 9092 35624 9104
rect 34664 9064 35624 9092
rect 34664 9052 34670 9064
rect 35618 9052 35624 9064
rect 35676 9052 35682 9104
rect 23569 9027 23627 9033
rect 23569 9024 23581 9027
rect 20640 8996 23581 9024
rect 23569 8993 23581 8996
rect 23615 8993 23627 9027
rect 23569 8987 23627 8993
rect 23658 8984 23664 9036
rect 23716 9024 23722 9036
rect 24581 9027 24639 9033
rect 24581 9024 24593 9027
rect 23716 8996 24593 9024
rect 23716 8984 23722 8996
rect 24581 8993 24593 8996
rect 24627 8993 24639 9027
rect 24581 8987 24639 8993
rect 26418 8984 26424 9036
rect 26476 8984 26482 9036
rect 26602 8984 26608 9036
rect 26660 9024 26666 9036
rect 27525 9027 27583 9033
rect 27525 9024 27537 9027
rect 26660 8996 27537 9024
rect 26660 8984 26666 8996
rect 27525 8993 27537 8996
rect 27571 8993 27583 9027
rect 27525 8987 27583 8993
rect 28534 8984 28540 9036
rect 28592 9024 28598 9036
rect 28592 8996 29700 9024
rect 28592 8984 28598 8996
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19260 8928 19441 8956
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19522 8959 19580 8965
rect 19522 8925 19534 8959
rect 19568 8925 19580 8959
rect 19522 8919 19580 8925
rect 19702 8916 19708 8968
rect 19760 8916 19766 8968
rect 19978 8965 19984 8968
rect 19935 8959 19984 8965
rect 19935 8925 19947 8959
rect 19981 8925 19984 8959
rect 19935 8919 19984 8925
rect 19978 8916 19984 8919
rect 20036 8916 20042 8968
rect 21910 8916 21916 8968
rect 21968 8916 21974 8968
rect 23293 8959 23351 8965
rect 23293 8925 23305 8959
rect 23339 8956 23351 8959
rect 23474 8956 23480 8968
rect 23339 8928 23480 8956
rect 23339 8925 23351 8928
rect 23293 8919 23351 8925
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 26786 8916 26792 8968
rect 26844 8956 26850 8968
rect 27249 8959 27307 8965
rect 27249 8956 27261 8959
rect 26844 8928 27261 8956
rect 26844 8916 26850 8928
rect 27249 8925 27261 8928
rect 27295 8925 27307 8959
rect 29546 8956 29552 8968
rect 28658 8928 29552 8956
rect 27249 8919 27307 8925
rect 29546 8916 29552 8928
rect 29604 8916 29610 8968
rect 17494 8848 17500 8900
rect 17552 8848 17558 8900
rect 18598 8848 18604 8900
rect 18656 8848 18662 8900
rect 19797 8891 19855 8897
rect 19797 8857 19809 8891
rect 19843 8888 19855 8891
rect 19843 8860 20760 8888
rect 19843 8857 19855 8860
rect 19797 8851 19855 8857
rect 18690 8820 18696 8832
rect 17236 8792 18696 8820
rect 15344 8780 15350 8792
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 18877 8823 18935 8829
rect 18877 8789 18889 8823
rect 18923 8820 18935 8823
rect 19426 8820 19432 8832
rect 18923 8792 19432 8820
rect 18923 8789 18935 8792
rect 18877 8783 18935 8789
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 20073 8823 20131 8829
rect 20073 8789 20085 8823
rect 20119 8820 20131 8823
rect 20622 8820 20628 8832
rect 20119 8792 20628 8820
rect 20119 8789 20131 8792
rect 20073 8783 20131 8789
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20732 8820 20760 8860
rect 20806 8848 20812 8900
rect 20864 8848 20870 8900
rect 22833 8891 22891 8897
rect 22833 8857 22845 8891
rect 22879 8888 22891 8891
rect 24486 8888 24492 8900
rect 22879 8860 24492 8888
rect 22879 8857 22891 8860
rect 22833 8851 22891 8857
rect 24486 8848 24492 8860
rect 24544 8848 24550 8900
rect 24854 8848 24860 8900
rect 24912 8848 24918 8900
rect 29672 8888 29700 8996
rect 29914 8984 29920 9036
rect 29972 8984 29978 9036
rect 30006 8984 30012 9036
rect 30064 9024 30070 9036
rect 30745 9027 30803 9033
rect 30745 9024 30757 9027
rect 30064 8996 30757 9024
rect 30064 8984 30070 8996
rect 30745 8993 30757 8996
rect 30791 9024 30803 9027
rect 31754 9024 31760 9036
rect 30791 8996 31760 9024
rect 30791 8993 30803 8996
rect 30745 8987 30803 8993
rect 31754 8984 31760 8996
rect 31812 8984 31818 9036
rect 32766 8984 32772 9036
rect 32824 9024 32830 9036
rect 32824 8996 33916 9024
rect 32824 8984 32830 8996
rect 29733 8959 29791 8965
rect 29733 8925 29745 8959
rect 29779 8956 29791 8959
rect 29932 8956 29960 8984
rect 29779 8928 29960 8956
rect 30101 8959 30159 8965
rect 29779 8925 29791 8928
rect 29733 8919 29791 8925
rect 30101 8925 30113 8959
rect 30147 8956 30159 8959
rect 30282 8956 30288 8968
rect 30147 8928 30288 8956
rect 30147 8925 30159 8928
rect 30101 8919 30159 8925
rect 30282 8916 30288 8928
rect 30340 8916 30346 8968
rect 33505 8959 33563 8965
rect 33505 8925 33517 8959
rect 33551 8956 33563 8959
rect 33594 8956 33600 8968
rect 33551 8928 33600 8956
rect 33551 8925 33563 8928
rect 33505 8919 33563 8925
rect 33594 8916 33600 8928
rect 33652 8916 33658 8968
rect 33686 8916 33692 8968
rect 33744 8916 33750 8968
rect 33888 8965 33916 8996
rect 34882 8984 34888 9036
rect 34940 9024 34946 9036
rect 35158 9024 35164 9036
rect 34940 8996 35164 9024
rect 34940 8984 34946 8996
rect 35158 8984 35164 8996
rect 35216 8984 35222 9036
rect 35342 8984 35348 9036
rect 35400 8984 35406 9036
rect 35526 8984 35532 9036
rect 35584 8984 35590 9036
rect 35894 8984 35900 9036
rect 35952 9024 35958 9036
rect 36817 9027 36875 9033
rect 36817 9024 36829 9027
rect 35952 8996 36829 9024
rect 35952 8984 35958 8996
rect 36817 8993 36829 8996
rect 36863 8993 36875 9027
rect 36817 8987 36875 8993
rect 33873 8959 33931 8965
rect 33873 8925 33885 8959
rect 33919 8925 33931 8959
rect 33873 8919 33931 8925
rect 35250 8916 35256 8968
rect 35308 8916 35314 8968
rect 35618 8916 35624 8968
rect 35676 8956 35682 8968
rect 36081 8959 36139 8965
rect 36081 8956 36093 8959
rect 35676 8928 36093 8956
rect 35676 8916 35682 8928
rect 36081 8925 36093 8928
rect 36127 8925 36139 8959
rect 36081 8919 36139 8925
rect 29914 8888 29920 8900
rect 26082 8860 27200 8888
rect 29672 8860 29920 8888
rect 22281 8823 22339 8829
rect 22281 8820 22293 8823
rect 20732 8792 22293 8820
rect 22281 8789 22293 8792
rect 22327 8820 22339 8823
rect 22462 8820 22468 8832
rect 22327 8792 22468 8820
rect 22327 8789 22339 8792
rect 22281 8783 22339 8789
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 23385 8823 23443 8829
rect 23385 8789 23397 8823
rect 23431 8820 23443 8823
rect 26418 8820 26424 8832
rect 23431 8792 26424 8820
rect 23431 8789 23443 8792
rect 23385 8783 23443 8789
rect 26418 8780 26424 8792
rect 26476 8780 26482 8832
rect 27172 8820 27200 8860
rect 29914 8848 29920 8860
rect 29972 8848 29978 8900
rect 30009 8891 30067 8897
rect 30009 8857 30021 8891
rect 30055 8888 30067 8891
rect 30190 8888 30196 8900
rect 30055 8860 30196 8888
rect 30055 8857 30067 8860
rect 30009 8851 30067 8857
rect 30190 8848 30196 8860
rect 30248 8848 30254 8900
rect 30466 8848 30472 8900
rect 30524 8888 30530 8900
rect 31021 8891 31079 8897
rect 31021 8888 31033 8891
rect 30524 8860 31033 8888
rect 30524 8848 30530 8860
rect 31021 8857 31033 8860
rect 31067 8857 31079 8891
rect 32246 8860 33732 8888
rect 31021 8851 31079 8857
rect 28902 8820 28908 8832
rect 27172 8792 28908 8820
rect 28902 8780 28908 8792
rect 28960 8780 28966 8832
rect 30742 8780 30748 8832
rect 30800 8820 30806 8832
rect 32493 8823 32551 8829
rect 32493 8820 32505 8823
rect 30800 8792 32505 8820
rect 30800 8780 30806 8792
rect 32493 8789 32505 8792
rect 32539 8789 32551 8823
rect 33704 8820 33732 8860
rect 33778 8848 33784 8900
rect 33836 8848 33842 8900
rect 33980 8860 34836 8888
rect 33980 8820 34008 8860
rect 33704 8792 34008 8820
rect 32493 8783 32551 8789
rect 34054 8780 34060 8832
rect 34112 8780 34118 8832
rect 34808 8820 34836 8860
rect 34882 8848 34888 8900
rect 34940 8888 34946 8900
rect 36722 8888 36728 8900
rect 34940 8860 36728 8888
rect 34940 8848 34946 8860
rect 36722 8848 36728 8860
rect 36780 8848 36786 8900
rect 37090 8848 37096 8900
rect 37148 8848 37154 8900
rect 37550 8848 37556 8900
rect 37608 8848 37614 8900
rect 35618 8820 35624 8832
rect 34808 8792 35624 8820
rect 35618 8780 35624 8792
rect 35676 8780 35682 8832
rect 1104 8730 39352 8752
rect 1104 8678 10472 8730
rect 10524 8678 10536 8730
rect 10588 8678 10600 8730
rect 10652 8678 10664 8730
rect 10716 8678 10728 8730
rect 10780 8678 19994 8730
rect 20046 8678 20058 8730
rect 20110 8678 20122 8730
rect 20174 8678 20186 8730
rect 20238 8678 20250 8730
rect 20302 8678 29516 8730
rect 29568 8678 29580 8730
rect 29632 8678 29644 8730
rect 29696 8678 29708 8730
rect 29760 8678 29772 8730
rect 29824 8678 39038 8730
rect 39090 8678 39102 8730
rect 39154 8678 39166 8730
rect 39218 8678 39230 8730
rect 39282 8678 39294 8730
rect 39346 8678 39352 8730
rect 1104 8656 39352 8678
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8585 2927 8619
rect 2869 8579 2927 8585
rect 3237 8619 3295 8625
rect 3237 8585 3249 8619
rect 3283 8616 3295 8619
rect 3326 8616 3332 8628
rect 3283 8588 3332 8616
rect 3283 8585 3295 8588
rect 3237 8579 3295 8585
rect 2884 8548 2912 8579
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 6270 8616 6276 8628
rect 4304 8588 6276 8616
rect 4304 8576 4310 8588
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 8938 8616 8944 8628
rect 6880 8588 8944 8616
rect 6880 8576 6886 8588
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 9548 8588 10364 8616
rect 9548 8576 9554 8588
rect 4525 8551 4583 8557
rect 4525 8548 4537 8551
rect 2884 8520 4537 8548
rect 4525 8517 4537 8520
rect 4571 8517 4583 8551
rect 4525 8511 4583 8517
rect 4614 8508 4620 8560
rect 4672 8548 4678 8560
rect 7009 8551 7067 8557
rect 4672 8520 5014 8548
rect 4672 8508 4678 8520
rect 7009 8517 7021 8551
rect 7055 8548 7067 8551
rect 7466 8548 7472 8560
rect 7055 8520 7472 8548
rect 7055 8517 7067 8520
rect 7009 8511 7067 8517
rect 7466 8508 7472 8520
rect 7524 8508 7530 8560
rect 8570 8508 8576 8560
rect 8628 8508 8634 8560
rect 10134 8548 10140 8560
rect 9798 8520 10140 8548
rect 10134 8508 10140 8520
rect 10192 8508 10198 8560
rect 10336 8557 10364 8588
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 11480 8588 12020 8616
rect 11480 8576 11486 8588
rect 10321 8551 10379 8557
rect 10321 8517 10333 8551
rect 10367 8517 10379 8551
rect 10321 8511 10379 8517
rect 10778 8508 10784 8560
rect 10836 8508 10842 8560
rect 10997 8551 11055 8557
rect 10997 8517 11009 8551
rect 11043 8548 11055 8551
rect 11043 8520 11836 8548
rect 11043 8517 11055 8520
rect 10997 8511 11055 8517
rect 934 8440 940 8492
rect 992 8480 998 8492
rect 1581 8483 1639 8489
rect 1581 8480 1593 8483
rect 992 8452 1593 8480
rect 992 8440 998 8452
rect 1581 8449 1593 8452
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2774 8480 2780 8492
rect 1903 8452 2780 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2774 8440 2780 8452
rect 2832 8480 2838 8492
rect 3142 8480 3148 8492
rect 2832 8452 3148 8480
rect 2832 8440 2838 8452
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8480 3387 8483
rect 3375 8452 4016 8480
rect 3375 8449 3387 8452
rect 3329 8443 3387 8449
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 3344 8412 3372 8443
rect 2004 8384 3372 8412
rect 2004 8372 2010 8384
rect 3418 8372 3424 8424
rect 3476 8372 3482 8424
rect 3988 8412 4016 8452
rect 4246 8440 4252 8492
rect 4304 8440 4310 8492
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6880 8452 6929 8480
rect 6880 8440 6886 8452
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 7926 8480 7932 8492
rect 7432 8452 7932 8480
rect 7432 8440 7438 8452
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11422 8480 11428 8492
rect 11296 8452 11428 8480
rect 11296 8440 11302 8452
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 5997 8415 6055 8421
rect 5997 8412 6009 8415
rect 3988 8384 6009 8412
rect 5997 8381 6009 8384
rect 6043 8381 6055 8415
rect 5997 8375 6055 8381
rect 6564 8384 7052 8412
rect 6564 8353 6592 8384
rect 6549 8347 6607 8353
rect 6549 8313 6561 8347
rect 6595 8313 6607 8347
rect 7024 8344 7052 8384
rect 7098 8372 7104 8424
rect 7156 8372 7162 8424
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 8110 8412 8116 8424
rect 7248 8384 8116 8412
rect 7248 8372 7254 8384
rect 8110 8372 8116 8384
rect 8168 8412 8174 8424
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 8168 8384 8309 8412
rect 8168 8372 8174 8384
rect 8297 8381 8309 8384
rect 8343 8381 8355 8415
rect 9766 8412 9772 8424
rect 8297 8375 8355 8381
rect 8404 8384 9772 8412
rect 8404 8344 8432 8384
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8381 11759 8415
rect 11808 8412 11836 8520
rect 11882 8440 11888 8492
rect 11940 8440 11946 8492
rect 11992 8480 12020 8588
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 12584 8588 13308 8616
rect 12584 8576 12590 8588
rect 12066 8508 12072 8560
rect 12124 8548 12130 8560
rect 12124 8520 12480 8548
rect 12124 8508 12130 8520
rect 12452 8489 12480 8520
rect 13170 8508 13176 8560
rect 13228 8508 13234 8560
rect 13280 8548 13308 8588
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14093 8619 14151 8625
rect 14093 8616 14105 8619
rect 13964 8588 14105 8616
rect 13964 8576 13970 8588
rect 14093 8585 14105 8588
rect 14139 8585 14151 8619
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14093 8579 14151 8585
rect 14200 8588 14565 8616
rect 14200 8548 14228 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14553 8579 14611 8585
rect 14918 8576 14924 8628
rect 14976 8616 14982 8628
rect 15378 8616 15384 8628
rect 14976 8588 15384 8616
rect 14976 8576 14982 8588
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 20717 8619 20775 8625
rect 20717 8616 20729 8619
rect 15804 8588 20729 8616
rect 15804 8576 15810 8588
rect 20717 8585 20729 8588
rect 20763 8585 20775 8619
rect 20717 8579 20775 8585
rect 20806 8576 20812 8628
rect 20864 8616 20870 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 20864 8588 22017 8616
rect 20864 8576 20870 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 22186 8576 22192 8628
rect 22244 8616 22250 8628
rect 22373 8619 22431 8625
rect 22373 8616 22385 8619
rect 22244 8588 22385 8616
rect 22244 8576 22250 8588
rect 22373 8585 22385 8588
rect 22419 8585 22431 8619
rect 22373 8579 22431 8585
rect 22462 8576 22468 8628
rect 22520 8576 22526 8628
rect 23569 8619 23627 8625
rect 23569 8585 23581 8619
rect 23615 8616 23627 8619
rect 23842 8616 23848 8628
rect 23615 8588 23848 8616
rect 23615 8585 23627 8588
rect 23569 8579 23627 8585
rect 23842 8576 23848 8588
rect 23900 8616 23906 8628
rect 23900 8588 24716 8616
rect 23900 8576 23906 8588
rect 13280 8520 14228 8548
rect 14274 8508 14280 8560
rect 14332 8548 14338 8560
rect 14461 8551 14519 8557
rect 14461 8548 14473 8551
rect 14332 8520 14473 8548
rect 14332 8508 14338 8520
rect 14461 8517 14473 8520
rect 14507 8548 14519 8551
rect 17034 8548 17040 8560
rect 14507 8520 17040 8548
rect 14507 8517 14519 8520
rect 14461 8511 14519 8517
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 17126 8508 17132 8560
rect 17184 8508 17190 8560
rect 17586 8508 17592 8560
rect 17644 8508 17650 8560
rect 24026 8548 24032 8560
rect 19306 8520 24032 8548
rect 12253 8483 12311 8489
rect 12253 8480 12265 8483
rect 11992 8452 12265 8480
rect 12253 8449 12265 8452
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 12713 8483 12771 8489
rect 12713 8480 12725 8483
rect 12676 8452 12725 8480
rect 12676 8440 12682 8452
rect 12713 8449 12725 8452
rect 12759 8480 12771 8483
rect 14826 8480 14832 8492
rect 12759 8452 14832 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15746 8480 15752 8492
rect 15304 8452 15752 8480
rect 13170 8412 13176 8424
rect 11808 8384 13176 8412
rect 11701 8375 11759 8381
rect 11149 8347 11207 8353
rect 7024 8316 8432 8344
rect 9646 8316 11100 8344
rect 6549 8307 6607 8313
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 5626 8276 5632 8288
rect 3384 8248 5632 8276
rect 3384 8236 3390 8248
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 9646 8276 9674 8316
rect 6880 8248 9674 8276
rect 6880 8236 6886 8248
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10778 8276 10784 8288
rect 10008 8248 10784 8276
rect 10008 8236 10014 8248
rect 10778 8236 10784 8248
rect 10836 8276 10842 8288
rect 10965 8279 11023 8285
rect 10965 8276 10977 8279
rect 10836 8248 10977 8276
rect 10836 8236 10842 8248
rect 10965 8245 10977 8248
rect 11011 8245 11023 8279
rect 11072 8276 11100 8316
rect 11149 8313 11161 8347
rect 11195 8344 11207 8347
rect 11716 8344 11744 8375
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 14608 8384 14657 8412
rect 14608 8372 14614 8384
rect 14645 8381 14657 8384
rect 14691 8381 14703 8415
rect 15304 8412 15332 8452
rect 15746 8440 15752 8452
rect 15804 8480 15810 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15804 8452 15945 8480
rect 15804 8440 15810 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 16025 8483 16083 8489
rect 16025 8449 16037 8483
rect 16071 8480 16083 8483
rect 16666 8480 16672 8492
rect 16071 8452 16672 8480
rect 16071 8449 16083 8452
rect 16025 8443 16083 8449
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16816 8452 16865 8480
rect 16816 8440 16822 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 14645 8375 14703 8381
rect 15212 8384 15332 8412
rect 14274 8344 14280 8356
rect 11195 8316 11744 8344
rect 13188 8316 14280 8344
rect 11195 8313 11207 8316
rect 11149 8307 11207 8313
rect 13188 8276 13216 8316
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 11072 8248 13216 8276
rect 10965 8239 11023 8245
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 15212 8276 15240 8384
rect 15378 8372 15384 8424
rect 15436 8412 15442 8424
rect 16209 8415 16267 8421
rect 16209 8412 16221 8415
rect 15436 8384 16221 8412
rect 15436 8372 15442 8384
rect 16209 8381 16221 8384
rect 16255 8412 16267 8415
rect 16390 8412 16396 8424
rect 16255 8384 16396 8412
rect 16255 8381 16267 8384
rect 16209 8375 16267 8381
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 19306 8412 19334 8520
rect 24026 8508 24032 8520
rect 24084 8508 24090 8560
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8480 19763 8483
rect 20346 8480 20352 8492
rect 19751 8452 20352 8480
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 21542 8440 21548 8492
rect 21600 8480 21606 8492
rect 23293 8483 23351 8489
rect 21600 8452 23152 8480
rect 21600 8440 21606 8452
rect 16592 8384 19334 8412
rect 19797 8415 19855 8421
rect 15565 8347 15623 8353
rect 15565 8313 15577 8347
rect 15611 8313 15623 8347
rect 15565 8307 15623 8313
rect 13320 8248 15240 8276
rect 15580 8276 15608 8307
rect 15746 8304 15752 8356
rect 15804 8344 15810 8356
rect 16022 8344 16028 8356
rect 15804 8316 16028 8344
rect 15804 8304 15810 8316
rect 16022 8304 16028 8316
rect 16080 8304 16086 8356
rect 16592 8276 16620 8384
rect 19797 8381 19809 8415
rect 19843 8381 19855 8415
rect 19797 8375 19855 8381
rect 18506 8304 18512 8356
rect 18564 8344 18570 8356
rect 19337 8347 19395 8353
rect 19337 8344 19349 8347
rect 18564 8316 19349 8344
rect 18564 8304 18570 8316
rect 19337 8313 19349 8316
rect 19383 8313 19395 8347
rect 19337 8307 19395 8313
rect 19426 8304 19432 8356
rect 19484 8344 19490 8356
rect 19812 8344 19840 8375
rect 19886 8372 19892 8424
rect 19944 8412 19950 8424
rect 19981 8415 20039 8421
rect 19981 8412 19993 8415
rect 19944 8384 19993 8412
rect 19944 8372 19950 8384
rect 19981 8381 19993 8384
rect 20027 8412 20039 8415
rect 20530 8412 20536 8424
rect 20027 8384 20536 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 20990 8372 20996 8424
rect 21048 8412 21054 8424
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 21048 8384 21189 8412
rect 21048 8372 21054 8384
rect 21177 8381 21189 8384
rect 21223 8381 21235 8415
rect 21177 8375 21235 8381
rect 21361 8415 21419 8421
rect 21361 8381 21373 8415
rect 21407 8412 21419 8415
rect 22649 8415 22707 8421
rect 22649 8412 22661 8415
rect 21407 8384 22661 8412
rect 21407 8381 21419 8384
rect 21361 8375 21419 8381
rect 22649 8381 22661 8384
rect 22695 8412 22707 8415
rect 23014 8412 23020 8424
rect 22695 8384 23020 8412
rect 22695 8381 22707 8384
rect 22649 8375 22707 8381
rect 23014 8372 23020 8384
rect 23072 8372 23078 8424
rect 23124 8412 23152 8452
rect 23293 8449 23305 8483
rect 23339 8480 23351 8483
rect 24394 8480 24400 8492
rect 23339 8452 24400 8480
rect 23339 8449 23351 8452
rect 23293 8443 23351 8449
rect 24394 8440 24400 8452
rect 24452 8440 24458 8492
rect 24688 8489 24716 8588
rect 24854 8576 24860 8628
rect 24912 8616 24918 8628
rect 25777 8619 25835 8625
rect 25777 8616 25789 8619
rect 24912 8588 25789 8616
rect 24912 8576 24918 8588
rect 25777 8585 25789 8588
rect 25823 8585 25835 8619
rect 25777 8579 25835 8585
rect 25958 8576 25964 8628
rect 26016 8616 26022 8628
rect 26145 8619 26203 8625
rect 26145 8616 26157 8619
rect 26016 8588 26157 8616
rect 26016 8576 26022 8588
rect 26145 8585 26157 8588
rect 26191 8585 26203 8619
rect 26145 8579 26203 8585
rect 26234 8576 26240 8628
rect 26292 8576 26298 8628
rect 26344 8588 28764 8616
rect 24762 8508 24768 8560
rect 24820 8548 24826 8560
rect 26344 8548 26372 8588
rect 24820 8520 26372 8548
rect 24820 8508 24826 8520
rect 27430 8508 27436 8560
rect 27488 8508 27494 8560
rect 28442 8508 28448 8560
rect 28500 8508 28506 8560
rect 28736 8548 28764 8588
rect 28902 8576 28908 8628
rect 28960 8576 28966 8628
rect 28994 8576 29000 8628
rect 29052 8616 29058 8628
rect 29822 8616 29828 8628
rect 29052 8588 29828 8616
rect 29052 8576 29058 8588
rect 29822 8576 29828 8588
rect 29880 8576 29886 8628
rect 29914 8576 29920 8628
rect 29972 8616 29978 8628
rect 31846 8616 31852 8628
rect 29972 8588 31852 8616
rect 29972 8576 29978 8588
rect 31846 8576 31852 8588
rect 31904 8576 31910 8628
rect 32306 8576 32312 8628
rect 32364 8576 32370 8628
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 32769 8619 32827 8625
rect 32769 8616 32781 8619
rect 32548 8588 32781 8616
rect 32548 8576 32554 8588
rect 32769 8585 32781 8588
rect 32815 8585 32827 8619
rect 32769 8579 32827 8585
rect 32858 8576 32864 8628
rect 32916 8616 32922 8628
rect 33410 8616 33416 8628
rect 32916 8588 33416 8616
rect 32916 8576 32922 8588
rect 33410 8576 33416 8588
rect 33468 8616 33474 8628
rect 33965 8619 34023 8625
rect 33965 8616 33977 8619
rect 33468 8588 33977 8616
rect 33468 8576 33474 8588
rect 33965 8585 33977 8588
rect 34011 8585 34023 8619
rect 33965 8579 34023 8585
rect 34698 8576 34704 8628
rect 34756 8616 34762 8628
rect 37461 8619 37519 8625
rect 37461 8616 37473 8619
rect 34756 8588 37473 8616
rect 34756 8576 34762 8588
rect 37461 8585 37473 8588
rect 37507 8585 37519 8619
rect 37461 8579 37519 8585
rect 37918 8576 37924 8628
rect 37976 8576 37982 8628
rect 30190 8548 30196 8560
rect 28736 8520 30196 8548
rect 30190 8508 30196 8520
rect 30248 8508 30254 8560
rect 31018 8508 31024 8560
rect 31076 8508 31082 8560
rect 31386 8508 31392 8560
rect 31444 8548 31450 8560
rect 31662 8548 31668 8560
rect 31444 8520 31668 8548
rect 31444 8508 31450 8520
rect 31662 8508 31668 8520
rect 31720 8508 31726 8560
rect 32677 8551 32735 8557
rect 32677 8517 32689 8551
rect 32723 8548 32735 8551
rect 33594 8548 33600 8560
rect 32723 8520 33600 8548
rect 32723 8517 32735 8520
rect 32677 8511 32735 8517
rect 33594 8508 33600 8520
rect 33652 8508 33658 8560
rect 33796 8520 35388 8548
rect 24673 8483 24731 8489
rect 24673 8449 24685 8483
rect 24719 8449 24731 8483
rect 24673 8443 24731 8449
rect 25225 8483 25283 8489
rect 25225 8449 25237 8483
rect 25271 8480 25283 8483
rect 25774 8480 25780 8492
rect 25271 8452 25780 8480
rect 25271 8449 25283 8452
rect 25225 8443 25283 8449
rect 25774 8440 25780 8452
rect 25832 8440 25838 8492
rect 28902 8440 28908 8492
rect 28960 8480 28966 8492
rect 29825 8483 29883 8489
rect 29825 8480 29837 8483
rect 28960 8452 29837 8480
rect 28960 8440 28966 8452
rect 29825 8449 29837 8452
rect 29871 8449 29883 8483
rect 29825 8443 29883 8449
rect 31113 8483 31171 8489
rect 31113 8449 31125 8483
rect 31159 8480 31171 8483
rect 33318 8480 33324 8492
rect 31159 8452 33324 8480
rect 31159 8449 31171 8452
rect 31113 8443 31171 8449
rect 33318 8440 33324 8452
rect 33376 8440 33382 8492
rect 25590 8412 25596 8424
rect 23124 8384 25596 8412
rect 25590 8372 25596 8384
rect 25648 8372 25654 8424
rect 26421 8415 26479 8421
rect 26421 8381 26433 8415
rect 26467 8412 26479 8415
rect 26510 8412 26516 8424
rect 26467 8384 26516 8412
rect 26467 8381 26479 8384
rect 26421 8375 26479 8381
rect 26510 8372 26516 8384
rect 26568 8372 26574 8424
rect 26786 8372 26792 8424
rect 26844 8412 26850 8424
rect 27157 8415 27215 8421
rect 27157 8412 27169 8415
rect 26844 8384 27169 8412
rect 26844 8372 26850 8384
rect 27157 8381 27169 8384
rect 27203 8381 27215 8415
rect 27890 8412 27896 8424
rect 27157 8375 27215 8381
rect 27264 8384 27896 8412
rect 19484 8316 19748 8344
rect 19812 8316 19937 8344
rect 19484 8304 19490 8316
rect 15580 8248 16620 8276
rect 13320 8236 13326 8248
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 17494 8276 17500 8288
rect 16724 8248 17500 8276
rect 16724 8236 16730 8248
rect 17494 8236 17500 8248
rect 17552 8276 17558 8288
rect 19610 8276 19616 8288
rect 17552 8248 19616 8276
rect 17552 8236 17558 8248
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 19720 8276 19748 8316
rect 19794 8276 19800 8288
rect 19720 8248 19800 8276
rect 19794 8236 19800 8248
rect 19852 8236 19858 8288
rect 19909 8276 19937 8316
rect 20254 8304 20260 8356
rect 20312 8344 20318 8356
rect 25498 8344 25504 8356
rect 20312 8316 25504 8344
rect 20312 8304 20318 8316
rect 25498 8304 25504 8316
rect 25556 8304 25562 8356
rect 25682 8304 25688 8356
rect 25740 8304 25746 8356
rect 25958 8304 25964 8356
rect 26016 8344 26022 8356
rect 27264 8344 27292 8384
rect 27890 8372 27896 8384
rect 27948 8412 27954 8424
rect 29917 8415 29975 8421
rect 29917 8412 29929 8415
rect 27948 8384 29929 8412
rect 27948 8372 27954 8384
rect 29917 8381 29929 8384
rect 29963 8381 29975 8415
rect 29917 8375 29975 8381
rect 30101 8415 30159 8421
rect 30101 8381 30113 8415
rect 30147 8412 30159 8415
rect 30282 8412 30288 8424
rect 30147 8384 30288 8412
rect 30147 8381 30159 8384
rect 30101 8375 30159 8381
rect 30282 8372 30288 8384
rect 30340 8372 30346 8424
rect 31202 8372 31208 8424
rect 31260 8372 31266 8424
rect 32950 8372 32956 8424
rect 33008 8372 33014 8424
rect 33796 8412 33824 8520
rect 33870 8440 33876 8492
rect 33928 8440 33934 8492
rect 34882 8440 34888 8492
rect 34940 8440 34946 8492
rect 35360 8480 35388 8520
rect 35434 8508 35440 8560
rect 35492 8548 35498 8560
rect 35492 8520 36216 8548
rect 35492 8508 35498 8520
rect 35360 8452 35940 8480
rect 33336 8384 33824 8412
rect 26016 8316 27292 8344
rect 26016 8304 26022 8316
rect 28810 8304 28816 8356
rect 28868 8344 28874 8356
rect 28994 8344 29000 8356
rect 28868 8316 29000 8344
rect 28868 8304 28874 8316
rect 28994 8304 29000 8316
rect 29052 8304 29058 8356
rect 29086 8304 29092 8356
rect 29144 8344 29150 8356
rect 29457 8347 29515 8353
rect 29457 8344 29469 8347
rect 29144 8316 29469 8344
rect 29144 8304 29150 8316
rect 29457 8313 29469 8316
rect 29503 8313 29515 8347
rect 29457 8307 29515 8313
rect 29546 8304 29552 8356
rect 29604 8344 29610 8356
rect 33336 8344 33364 8384
rect 34054 8372 34060 8424
rect 34112 8372 34118 8424
rect 35158 8372 35164 8424
rect 35216 8412 35222 8424
rect 35526 8412 35532 8424
rect 35216 8384 35532 8412
rect 35216 8372 35222 8384
rect 35526 8372 35532 8384
rect 35584 8372 35590 8424
rect 35912 8412 35940 8452
rect 35986 8440 35992 8492
rect 36044 8440 36050 8492
rect 36188 8489 36216 8520
rect 36173 8483 36231 8489
rect 36173 8449 36185 8483
rect 36219 8449 36231 8483
rect 36173 8443 36231 8449
rect 37826 8440 37832 8492
rect 37884 8440 37890 8492
rect 36906 8412 36912 8424
rect 35912 8384 36912 8412
rect 36906 8372 36912 8384
rect 36964 8372 36970 8424
rect 38013 8415 38071 8421
rect 38013 8381 38025 8415
rect 38059 8381 38071 8415
rect 38013 8375 38071 8381
rect 29604 8316 33364 8344
rect 29604 8304 29610 8316
rect 33410 8304 33416 8356
rect 33468 8344 33474 8356
rect 33505 8347 33563 8353
rect 33505 8344 33517 8347
rect 33468 8316 33517 8344
rect 33468 8304 33474 8316
rect 33505 8313 33517 8316
rect 33551 8313 33563 8347
rect 33505 8307 33563 8313
rect 33612 8316 35296 8344
rect 21450 8276 21456 8288
rect 19909 8248 21456 8276
rect 21450 8236 21456 8248
rect 21508 8236 21514 8288
rect 25130 8236 25136 8288
rect 25188 8276 25194 8288
rect 25700 8276 25728 8304
rect 30190 8276 30196 8288
rect 25188 8248 30196 8276
rect 25188 8236 25194 8248
rect 30190 8236 30196 8248
rect 30248 8236 30254 8288
rect 30653 8279 30711 8285
rect 30653 8245 30665 8279
rect 30699 8276 30711 8279
rect 31662 8276 31668 8288
rect 30699 8248 31668 8276
rect 30699 8245 30711 8248
rect 30653 8239 30711 8245
rect 31662 8236 31668 8248
rect 31720 8236 31726 8288
rect 33042 8236 33048 8288
rect 33100 8276 33106 8288
rect 33612 8276 33640 8316
rect 33100 8248 33640 8276
rect 33100 8236 33106 8248
rect 33778 8236 33784 8288
rect 33836 8276 33842 8288
rect 34054 8276 34060 8288
rect 33836 8248 34060 8276
rect 33836 8236 33842 8248
rect 34054 8236 34060 8248
rect 34112 8236 34118 8288
rect 34882 8236 34888 8288
rect 34940 8276 34946 8288
rect 35158 8276 35164 8288
rect 34940 8248 35164 8276
rect 34940 8236 34946 8248
rect 35158 8236 35164 8248
rect 35216 8236 35222 8288
rect 35268 8276 35296 8316
rect 35342 8304 35348 8356
rect 35400 8344 35406 8356
rect 36357 8347 36415 8353
rect 36357 8344 36369 8347
rect 35400 8316 36369 8344
rect 35400 8304 35406 8316
rect 36357 8313 36369 8316
rect 36403 8313 36415 8347
rect 38028 8344 38056 8375
rect 36357 8307 36415 8313
rect 36464 8316 38056 8344
rect 36464 8276 36492 8316
rect 35268 8248 36492 8276
rect 1104 8186 39192 8208
rect 1104 8134 5711 8186
rect 5763 8134 5775 8186
rect 5827 8134 5839 8186
rect 5891 8134 5903 8186
rect 5955 8134 5967 8186
rect 6019 8134 15233 8186
rect 15285 8134 15297 8186
rect 15349 8134 15361 8186
rect 15413 8134 15425 8186
rect 15477 8134 15489 8186
rect 15541 8134 24755 8186
rect 24807 8134 24819 8186
rect 24871 8134 24883 8186
rect 24935 8134 24947 8186
rect 24999 8134 25011 8186
rect 25063 8134 34277 8186
rect 34329 8134 34341 8186
rect 34393 8134 34405 8186
rect 34457 8134 34469 8186
rect 34521 8134 34533 8186
rect 34585 8134 39192 8186
rect 1104 8112 39192 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2958 8072 2964 8084
rect 2179 8044 2964 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2958 8032 2964 8044
rect 3016 8072 3022 8084
rect 3016 8044 3280 8072
rect 3016 8032 3022 8044
rect 2317 8007 2375 8013
rect 2317 7973 2329 8007
rect 2363 8004 2375 8007
rect 3252 8004 3280 8044
rect 3326 8032 3332 8084
rect 3384 8072 3390 8084
rect 3973 8075 4031 8081
rect 3973 8072 3985 8075
rect 3384 8044 3985 8072
rect 3384 8032 3390 8044
rect 3973 8041 3985 8044
rect 4019 8041 4031 8075
rect 3973 8035 4031 8041
rect 4430 8032 4436 8084
rect 4488 8032 4494 8084
rect 9030 8072 9036 8084
rect 5552 8044 9036 8072
rect 3878 8004 3884 8016
rect 2363 7976 2774 8004
rect 3252 7976 3884 8004
rect 2363 7973 2375 7976
rect 2317 7967 2375 7973
rect 2746 7936 2774 7976
rect 3878 7964 3884 7976
rect 3936 7964 3942 8016
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 2746 7908 4077 7936
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4614 7936 4620 7948
rect 4065 7899 4123 7905
rect 4172 7908 4620 7936
rect 2774 7828 2780 7880
rect 2832 7828 2838 7880
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 4172 7868 4200 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 5552 7945 5580 8044
rect 9030 8032 9036 8044
rect 9088 8072 9094 8084
rect 9088 8044 9444 8072
rect 9088 8032 9094 8044
rect 5537 7939 5595 7945
rect 5537 7905 5549 7939
rect 5583 7905 5595 7939
rect 5537 7899 5595 7905
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 7098 7936 7104 7948
rect 6328 7908 7104 7936
rect 6328 7896 6334 7908
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 8846 7936 8852 7948
rect 7616 7908 8852 7936
rect 7616 7896 7622 7908
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 9416 7936 9444 8044
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 10836 8044 13461 8072
rect 10836 8032 10842 8044
rect 13449 8041 13461 8044
rect 13495 8072 13507 8075
rect 13495 8044 14320 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 12342 7964 12348 8016
rect 12400 8004 12406 8016
rect 13633 8007 13691 8013
rect 13633 8004 13645 8007
rect 12400 7976 13645 8004
rect 12400 7964 12406 7976
rect 13633 7973 13645 7976
rect 13679 7973 13691 8007
rect 14292 8004 14320 8044
rect 14366 8032 14372 8084
rect 14424 8032 14430 8084
rect 16298 8072 16304 8084
rect 14476 8044 16304 8072
rect 14476 8004 14504 8044
rect 16298 8032 16304 8044
rect 16356 8072 16362 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 16356 8044 17693 8072
rect 16356 8032 16362 8044
rect 17681 8041 17693 8044
rect 17727 8072 17739 8075
rect 17770 8072 17776 8084
rect 17727 8044 17776 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 17865 8075 17923 8081
rect 17865 8041 17877 8075
rect 17911 8072 17923 8075
rect 17954 8072 17960 8084
rect 17911 8044 17960 8072
rect 17911 8041 17923 8044
rect 17865 8035 17923 8041
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18877 8075 18935 8081
rect 18877 8072 18889 8075
rect 18196 8044 18889 8072
rect 18196 8032 18202 8044
rect 18877 8041 18889 8044
rect 18923 8041 18935 8075
rect 18877 8035 18935 8041
rect 18966 8032 18972 8084
rect 19024 8072 19030 8084
rect 19024 8044 22232 8072
rect 19024 8032 19030 8044
rect 14292 7976 14504 8004
rect 13633 7967 13691 7973
rect 14550 7964 14556 8016
rect 14608 8004 14614 8016
rect 15838 8004 15844 8016
rect 14608 7976 15844 8004
rect 14608 7964 14614 7976
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 19426 8004 19432 8016
rect 15948 7976 19432 8004
rect 9769 7939 9827 7945
rect 9769 7936 9781 7939
rect 9416 7908 9781 7936
rect 9769 7905 9781 7908
rect 9815 7936 9827 7939
rect 10686 7936 10692 7948
rect 9815 7908 10692 7936
rect 9815 7905 9827 7908
rect 9769 7899 9827 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 11054 7896 11060 7948
rect 11112 7896 11118 7948
rect 12802 7896 12808 7948
rect 12860 7896 12866 7948
rect 13648 7908 15148 7936
rect 13648 7880 13676 7908
rect 3896 7840 4200 7868
rect 4249 7871 4307 7877
rect 1946 7760 1952 7812
rect 2004 7760 2010 7812
rect 2130 7760 2136 7812
rect 2188 7809 2194 7812
rect 2188 7803 2223 7809
rect 2211 7800 2223 7803
rect 2682 7800 2688 7812
rect 2211 7772 2688 7800
rect 2211 7769 2223 7772
rect 2188 7763 2223 7769
rect 2188 7760 2194 7763
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 2961 7803 3019 7809
rect 2961 7769 2973 7803
rect 3007 7769 3019 7803
rect 2961 7763 3019 7769
rect 3053 7803 3111 7809
rect 3053 7769 3065 7803
rect 3099 7769 3111 7803
rect 3896 7800 3924 7840
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4338 7868 4344 7880
rect 4295 7840 4344 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5626 7868 5632 7880
rect 5307 7840 5632 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 9122 7868 9128 7880
rect 8628 7840 9128 7868
rect 8628 7828 8634 7840
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 3053 7763 3111 7769
rect 3252 7772 3924 7800
rect 3973 7803 4031 7809
rect 2406 7692 2412 7744
rect 2464 7732 2470 7744
rect 2976 7732 3004 7763
rect 2464 7704 3004 7732
rect 3068 7732 3096 7763
rect 3252 7732 3280 7772
rect 3973 7769 3985 7803
rect 4019 7800 4031 7803
rect 4706 7800 4712 7812
rect 4019 7772 4712 7800
rect 4019 7769 4031 7772
rect 3973 7763 4031 7769
rect 4706 7760 4712 7772
rect 4764 7760 4770 7812
rect 6549 7803 6607 7809
rect 6549 7800 6561 7803
rect 4908 7772 6561 7800
rect 3068 7704 3280 7732
rect 3329 7735 3387 7741
rect 2464 7692 2470 7704
rect 3329 7701 3341 7735
rect 3375 7732 3387 7735
rect 3878 7732 3884 7744
rect 3375 7704 3884 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4908 7741 4936 7772
rect 6549 7769 6561 7772
rect 6595 7769 6607 7803
rect 6549 7763 6607 7769
rect 7282 7760 7288 7812
rect 7340 7760 7346 7812
rect 8478 7760 8484 7812
rect 8536 7800 8542 7812
rect 9493 7803 9551 7809
rect 9493 7800 9505 7803
rect 8536 7772 9505 7800
rect 8536 7760 8542 7772
rect 9493 7769 9505 7772
rect 9539 7769 9551 7803
rect 10796 7800 10824 7831
rect 13630 7828 13636 7880
rect 13688 7828 13694 7880
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 14550 7868 14556 7880
rect 14323 7840 14556 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 14550 7828 14556 7840
rect 14608 7828 14614 7880
rect 14921 7871 14979 7877
rect 14921 7837 14933 7871
rect 14967 7868 14979 7871
rect 15010 7868 15016 7880
rect 14967 7840 15016 7868
rect 14967 7837 14979 7840
rect 14921 7831 14979 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15120 7868 15148 7908
rect 15194 7896 15200 7948
rect 15252 7936 15258 7948
rect 15562 7936 15568 7948
rect 15252 7908 15568 7936
rect 15252 7896 15258 7908
rect 15562 7896 15568 7908
rect 15620 7936 15626 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15620 7908 15669 7936
rect 15620 7896 15626 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 15948 7936 15976 7976
rect 19426 7964 19432 7976
rect 19484 7964 19490 8016
rect 22204 8004 22232 8044
rect 22278 8032 22284 8084
rect 22336 8072 22342 8084
rect 24581 8075 24639 8081
rect 22336 8044 23888 8072
rect 22336 8032 22342 8044
rect 23750 8004 23756 8016
rect 22204 7976 23756 8004
rect 23750 7964 23756 7976
rect 23808 7964 23814 8016
rect 15804 7908 15976 7936
rect 15804 7896 15810 7908
rect 16758 7896 16764 7948
rect 16816 7896 16822 7948
rect 16850 7896 16856 7948
rect 16908 7896 16914 7948
rect 23474 7936 23480 7948
rect 18340 7908 23480 7936
rect 15120 7840 17632 7868
rect 10962 7800 10968 7812
rect 10796 7772 10968 7800
rect 9493 7763 9551 7769
rect 10962 7760 10968 7772
rect 11020 7760 11026 7812
rect 11514 7760 11520 7812
rect 11572 7760 11578 7812
rect 13265 7803 13323 7809
rect 13265 7769 13277 7803
rect 13311 7800 13323 7803
rect 15746 7800 15752 7812
rect 13311 7772 15752 7800
rect 13311 7769 13323 7772
rect 13265 7763 13323 7769
rect 15746 7760 15752 7772
rect 15804 7760 15810 7812
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 16669 7803 16727 7809
rect 16669 7800 16681 7803
rect 16632 7772 16681 7800
rect 16632 7760 16638 7772
rect 16669 7769 16681 7772
rect 16715 7769 16727 7803
rect 16669 7763 16727 7769
rect 17494 7760 17500 7812
rect 17552 7760 17558 7812
rect 17604 7800 17632 7840
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 17954 7868 17960 7880
rect 17828 7840 17960 7868
rect 17828 7828 17834 7840
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18340 7877 18368 7908
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 23860 7945 23888 8044
rect 24581 8041 24593 8075
rect 24627 8072 24639 8075
rect 29990 8075 30048 8081
rect 29990 8072 30002 8075
rect 24627 8044 30002 8072
rect 24627 8041 24639 8044
rect 24581 8035 24639 8041
rect 29990 8041 30002 8044
rect 30036 8041 30048 8075
rect 29990 8035 30048 8041
rect 30190 8032 30196 8084
rect 30248 8072 30254 8084
rect 31481 8075 31539 8081
rect 31481 8072 31493 8075
rect 30248 8044 31493 8072
rect 30248 8032 30254 8044
rect 31481 8041 31493 8044
rect 31527 8041 31539 8075
rect 31481 8035 31539 8041
rect 32048 8044 33272 8072
rect 23934 7964 23940 8016
rect 23992 8004 23998 8016
rect 29086 8004 29092 8016
rect 23992 7976 25820 8004
rect 23992 7964 23998 7976
rect 23845 7939 23903 7945
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 24762 7936 24768 7948
rect 23891 7908 24768 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24762 7896 24768 7908
rect 24820 7896 24826 7948
rect 24854 7896 24860 7948
rect 24912 7936 24918 7948
rect 25225 7939 25283 7945
rect 25225 7936 25237 7939
rect 24912 7908 25237 7936
rect 24912 7896 24918 7908
rect 25225 7905 25237 7908
rect 25271 7936 25283 7939
rect 25271 7908 25728 7936
rect 25271 7905 25283 7908
rect 25225 7899 25283 7905
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18690 7828 18696 7880
rect 18748 7828 18754 7880
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19797 7871 19855 7877
rect 19797 7868 19809 7871
rect 19392 7840 19809 7868
rect 19392 7828 19398 7840
rect 19797 7837 19809 7840
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7868 22155 7871
rect 22186 7868 22192 7880
rect 22143 7840 22192 7868
rect 22143 7837 22155 7840
rect 22097 7831 22155 7837
rect 22186 7828 22192 7840
rect 22244 7828 22250 7880
rect 23290 7828 23296 7880
rect 23348 7868 23354 7880
rect 24946 7868 24952 7880
rect 23348 7840 24952 7868
rect 23348 7828 23354 7840
rect 24946 7828 24952 7840
rect 25004 7828 25010 7880
rect 18509 7803 18567 7809
rect 18509 7800 18521 7803
rect 17604 7772 18521 7800
rect 18509 7769 18521 7772
rect 18555 7769 18567 7803
rect 18509 7763 18567 7769
rect 18598 7760 18604 7812
rect 18656 7760 18662 7812
rect 18782 7760 18788 7812
rect 18840 7800 18846 7812
rect 20073 7803 20131 7809
rect 20073 7800 20085 7803
rect 18840 7772 20085 7800
rect 18840 7760 18846 7772
rect 20073 7769 20085 7772
rect 20119 7769 20131 7803
rect 20073 7763 20131 7769
rect 20714 7760 20720 7812
rect 20772 7760 20778 7812
rect 22465 7803 22523 7809
rect 22465 7800 22477 7803
rect 21376 7772 22477 7800
rect 4893 7735 4951 7741
rect 4893 7701 4905 7735
rect 4939 7701 4951 7735
rect 4893 7695 4951 7701
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 5353 7735 5411 7741
rect 5353 7732 5365 7735
rect 5132 7704 5365 7732
rect 5132 7692 5138 7704
rect 5353 7701 5365 7704
rect 5399 7732 5411 7735
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 5399 7704 8033 7732
rect 5399 7701 5411 7704
rect 5353 7695 5411 7701
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 9122 7692 9128 7744
rect 9180 7692 9186 7744
rect 9582 7692 9588 7744
rect 9640 7692 9646 7744
rect 13170 7692 13176 7744
rect 13228 7732 13234 7744
rect 13475 7735 13533 7741
rect 13475 7732 13487 7735
rect 13228 7704 13487 7732
rect 13228 7692 13234 7704
rect 13475 7701 13487 7704
rect 13521 7732 13533 7735
rect 14274 7732 14280 7744
rect 13521 7704 14280 7732
rect 13521 7701 13533 7704
rect 13475 7695 13533 7701
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 14458 7692 14464 7744
rect 14516 7732 14522 7744
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 14516 7704 16313 7732
rect 14516 7692 14522 7704
rect 16301 7701 16313 7704
rect 16347 7701 16359 7735
rect 16301 7695 16359 7701
rect 17707 7735 17765 7741
rect 17707 7701 17719 7735
rect 17753 7732 17765 7735
rect 17954 7732 17960 7744
rect 17753 7704 17960 7732
rect 17753 7701 17765 7704
rect 17707 7695 17765 7701
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 19610 7692 19616 7744
rect 19668 7732 19674 7744
rect 20254 7732 20260 7744
rect 19668 7704 20260 7732
rect 19668 7692 19674 7704
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 20438 7692 20444 7744
rect 20496 7732 20502 7744
rect 21376 7732 21404 7772
rect 22465 7769 22477 7772
rect 22511 7769 22523 7803
rect 22465 7763 22523 7769
rect 23569 7803 23627 7809
rect 23569 7769 23581 7803
rect 23615 7800 23627 7803
rect 23934 7800 23940 7812
rect 23615 7772 23940 7800
rect 23615 7769 23627 7772
rect 23569 7763 23627 7769
rect 23934 7760 23940 7772
rect 23992 7800 23998 7812
rect 24670 7800 24676 7812
rect 23992 7772 24676 7800
rect 23992 7760 23998 7772
rect 24670 7760 24676 7772
rect 24728 7760 24734 7812
rect 25041 7803 25099 7809
rect 25041 7769 25053 7803
rect 25087 7800 25099 7803
rect 25130 7800 25136 7812
rect 25087 7772 25136 7800
rect 25087 7769 25099 7772
rect 25041 7763 25099 7769
rect 25130 7760 25136 7772
rect 25188 7760 25194 7812
rect 25222 7760 25228 7812
rect 25280 7800 25286 7812
rect 25498 7800 25504 7812
rect 25280 7772 25504 7800
rect 25280 7760 25286 7772
rect 25498 7760 25504 7772
rect 25556 7760 25562 7812
rect 20496 7704 21404 7732
rect 20496 7692 20502 7704
rect 21542 7692 21548 7744
rect 21600 7692 21606 7744
rect 22646 7692 22652 7744
rect 22704 7732 22710 7744
rect 23201 7735 23259 7741
rect 23201 7732 23213 7735
rect 22704 7704 23213 7732
rect 22704 7692 22710 7704
rect 23201 7701 23213 7704
rect 23247 7701 23259 7735
rect 23201 7695 23259 7701
rect 23661 7735 23719 7741
rect 23661 7701 23673 7735
rect 23707 7732 23719 7735
rect 23842 7732 23848 7744
rect 23707 7704 23848 7732
rect 23707 7701 23719 7704
rect 23661 7695 23719 7701
rect 23842 7692 23848 7704
rect 23900 7692 23906 7744
rect 24949 7735 25007 7741
rect 24949 7701 24961 7735
rect 24995 7732 25007 7735
rect 25314 7732 25320 7744
rect 24995 7704 25320 7732
rect 24995 7701 25007 7704
rect 24949 7695 25007 7701
rect 25314 7692 25320 7704
rect 25372 7732 25378 7744
rect 25590 7732 25596 7744
rect 25372 7704 25596 7732
rect 25372 7692 25378 7704
rect 25590 7692 25596 7704
rect 25648 7692 25654 7744
rect 25700 7732 25728 7908
rect 25792 7877 25820 7976
rect 28276 7976 29092 8004
rect 26050 7896 26056 7948
rect 26108 7936 26114 7948
rect 26418 7936 26424 7948
rect 26108 7908 26424 7936
rect 26108 7896 26114 7908
rect 26418 7896 26424 7908
rect 26476 7896 26482 7948
rect 27065 7939 27123 7945
rect 27065 7905 27077 7939
rect 27111 7936 27123 7939
rect 28276 7936 28304 7976
rect 29086 7964 29092 7976
rect 29144 7964 29150 8016
rect 31386 7964 31392 8016
rect 31444 8004 31450 8016
rect 32048 8004 32076 8044
rect 31444 7976 32076 8004
rect 33244 8004 33272 8044
rect 33318 8032 33324 8084
rect 33376 8072 33382 8084
rect 33689 8075 33747 8081
rect 33689 8072 33701 8075
rect 33376 8044 33701 8072
rect 33376 8032 33382 8044
rect 33689 8041 33701 8044
rect 33735 8072 33747 8075
rect 34054 8072 34060 8084
rect 33735 8044 34060 8072
rect 33735 8041 33747 8044
rect 33689 8035 33747 8041
rect 34054 8032 34060 8044
rect 34112 8032 34118 8084
rect 34514 8032 34520 8084
rect 34572 8072 34578 8084
rect 35069 8075 35127 8081
rect 35069 8072 35081 8075
rect 34572 8044 35081 8072
rect 34572 8032 34578 8044
rect 35069 8041 35081 8044
rect 35115 8041 35127 8075
rect 35069 8035 35127 8041
rect 34146 8004 34152 8016
rect 33244 7976 34152 8004
rect 31444 7964 31450 7976
rect 34146 7964 34152 7976
rect 34204 8004 34210 8016
rect 35802 8004 35808 8016
rect 34204 7976 35808 8004
rect 34204 7964 34210 7976
rect 35802 7964 35808 7976
rect 35860 7964 35866 8016
rect 37734 7964 37740 8016
rect 37792 7964 37798 8016
rect 27111 7908 28304 7936
rect 28552 7908 28948 7936
rect 27111 7905 27123 7908
rect 27065 7899 27123 7905
rect 25777 7871 25835 7877
rect 25777 7837 25789 7871
rect 25823 7837 25835 7871
rect 25777 7831 25835 7837
rect 25866 7828 25872 7880
rect 25924 7868 25930 7880
rect 26145 7871 26203 7877
rect 26145 7868 26157 7871
rect 25924 7840 26157 7868
rect 25924 7828 25930 7840
rect 26145 7837 26157 7840
rect 26191 7868 26203 7871
rect 26602 7868 26608 7880
rect 26191 7840 26608 7868
rect 26191 7837 26203 7840
rect 26145 7831 26203 7837
rect 26602 7828 26608 7840
rect 26660 7828 26666 7880
rect 26786 7828 26792 7880
rect 26844 7828 26850 7880
rect 28552 7868 28580 7908
rect 28198 7840 28580 7868
rect 28810 7828 28816 7880
rect 28868 7828 28874 7880
rect 28920 7868 28948 7908
rect 28994 7896 29000 7948
rect 29052 7936 29058 7948
rect 29733 7939 29791 7945
rect 29733 7936 29745 7939
rect 29052 7908 29745 7936
rect 29052 7896 29058 7908
rect 29733 7905 29745 7908
rect 29779 7936 29791 7939
rect 30006 7936 30012 7948
rect 29779 7908 30012 7936
rect 29779 7905 29791 7908
rect 29733 7899 29791 7905
rect 30006 7896 30012 7908
rect 30064 7896 30070 7948
rect 31754 7896 31760 7948
rect 31812 7936 31818 7948
rect 31941 7939 31999 7945
rect 31941 7936 31953 7939
rect 31812 7908 31953 7936
rect 31812 7896 31818 7908
rect 31941 7905 31953 7908
rect 31987 7936 31999 7939
rect 33226 7936 33232 7948
rect 31987 7908 33232 7936
rect 31987 7905 31999 7908
rect 31941 7899 31999 7905
rect 33226 7896 33232 7908
rect 33284 7896 33290 7948
rect 33962 7896 33968 7948
rect 34020 7936 34026 7948
rect 34020 7908 35112 7936
rect 34020 7896 34026 7908
rect 34149 7871 34207 7877
rect 28920 7840 29776 7868
rect 25958 7760 25964 7812
rect 26016 7760 26022 7812
rect 26050 7760 26056 7812
rect 26108 7760 26114 7812
rect 26160 7772 26464 7800
rect 26160 7732 26188 7772
rect 25700 7704 26188 7732
rect 26326 7692 26332 7744
rect 26384 7692 26390 7744
rect 26436 7732 26464 7772
rect 28718 7732 28724 7744
rect 26436 7704 28724 7732
rect 28718 7692 28724 7704
rect 28776 7692 28782 7744
rect 28902 7692 28908 7744
rect 28960 7732 28966 7744
rect 29086 7732 29092 7744
rect 28960 7704 29092 7732
rect 28960 7692 28966 7704
rect 29086 7692 29092 7704
rect 29144 7692 29150 7744
rect 29748 7732 29776 7840
rect 33700 7840 34008 7868
rect 31234 7772 31616 7800
rect 31294 7732 31300 7744
rect 29748 7704 31300 7732
rect 31294 7692 31300 7704
rect 31352 7692 31358 7744
rect 31588 7732 31616 7772
rect 31662 7760 31668 7812
rect 31720 7800 31726 7812
rect 32217 7803 32275 7809
rect 32217 7800 32229 7803
rect 31720 7772 32229 7800
rect 31720 7760 31726 7772
rect 32217 7769 32229 7772
rect 32263 7769 32275 7803
rect 32217 7763 32275 7769
rect 32950 7760 32956 7812
rect 33008 7760 33014 7812
rect 33700 7732 33728 7840
rect 33980 7800 34008 7840
rect 34149 7837 34161 7871
rect 34195 7868 34207 7871
rect 34698 7868 34704 7880
rect 34195 7840 34704 7868
rect 34195 7837 34207 7840
rect 34149 7831 34207 7837
rect 34698 7828 34704 7840
rect 34756 7828 34762 7880
rect 35084 7877 35112 7908
rect 35158 7896 35164 7948
rect 35216 7896 35222 7948
rect 35894 7896 35900 7948
rect 35952 7936 35958 7948
rect 35989 7939 36047 7945
rect 35989 7936 36001 7939
rect 35952 7908 36001 7936
rect 35952 7896 35958 7908
rect 35989 7905 36001 7908
rect 36035 7905 36047 7939
rect 35989 7899 36047 7905
rect 35069 7871 35127 7877
rect 35069 7837 35081 7871
rect 35115 7837 35127 7871
rect 35069 7831 35127 7837
rect 35342 7828 35348 7880
rect 35400 7828 35406 7880
rect 34241 7803 34299 7809
rect 34241 7800 34253 7803
rect 33980 7772 34253 7800
rect 34241 7769 34253 7772
rect 34287 7769 34299 7803
rect 36004 7800 36032 7899
rect 36998 7896 37004 7948
rect 37056 7936 37062 7948
rect 37056 7908 38516 7936
rect 37056 7896 37062 7908
rect 37366 7828 37372 7880
rect 37424 7828 37430 7880
rect 38488 7877 38516 7908
rect 38473 7871 38531 7877
rect 38473 7837 38485 7871
rect 38519 7837 38531 7871
rect 38473 7831 38531 7837
rect 36170 7800 36176 7812
rect 36004 7772 36176 7800
rect 34241 7763 34299 7769
rect 36170 7760 36176 7772
rect 36228 7760 36234 7812
rect 36262 7760 36268 7812
rect 36320 7760 36326 7812
rect 38654 7760 38660 7812
rect 38712 7760 38718 7812
rect 31588 7704 33728 7732
rect 35526 7692 35532 7744
rect 35584 7692 35590 7744
rect 1104 7642 39352 7664
rect 1104 7590 10472 7642
rect 10524 7590 10536 7642
rect 10588 7590 10600 7642
rect 10652 7590 10664 7642
rect 10716 7590 10728 7642
rect 10780 7590 19994 7642
rect 20046 7590 20058 7642
rect 20110 7590 20122 7642
rect 20174 7590 20186 7642
rect 20238 7590 20250 7642
rect 20302 7590 29516 7642
rect 29568 7590 29580 7642
rect 29632 7590 29644 7642
rect 29696 7590 29708 7642
rect 29760 7590 29772 7642
rect 29824 7590 39038 7642
rect 39090 7590 39102 7642
rect 39154 7590 39166 7642
rect 39218 7590 39230 7642
rect 39282 7590 39294 7642
rect 39346 7590 39352 7642
rect 1104 7568 39352 7590
rect 3326 7488 3332 7540
rect 3384 7488 3390 7540
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 4798 7528 4804 7540
rect 4488 7500 4804 7528
rect 4488 7488 4494 7500
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 5629 7531 5687 7537
rect 5629 7497 5641 7531
rect 5675 7528 5687 7531
rect 7558 7528 7564 7540
rect 5675 7500 7564 7528
rect 5675 7497 5687 7500
rect 5629 7491 5687 7497
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 15010 7528 15016 7540
rect 7708 7500 15016 7528
rect 7708 7488 7714 7500
rect 2406 7420 2412 7472
rect 2464 7460 2470 7472
rect 2961 7463 3019 7469
rect 2961 7460 2973 7463
rect 2464 7432 2973 7460
rect 2464 7420 2470 7432
rect 2961 7429 2973 7432
rect 3007 7460 3019 7463
rect 3602 7460 3608 7472
rect 3007 7432 3608 7460
rect 3007 7429 3019 7432
rect 2961 7423 3019 7429
rect 3602 7420 3608 7432
rect 3660 7420 3666 7472
rect 6454 7460 6460 7472
rect 4080 7432 6460 7460
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 2041 7395 2099 7401
rect 2041 7392 2053 7395
rect 1728 7364 2053 7392
rect 1728 7352 1734 7364
rect 2041 7361 2053 7364
rect 2087 7361 2099 7395
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2041 7355 2099 7361
rect 2700 7364 2789 7392
rect 2222 7148 2228 7200
rect 2280 7148 2286 7200
rect 2700 7188 2728 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 3050 7352 3056 7404
rect 3108 7352 3114 7404
rect 3142 7352 3148 7404
rect 3200 7392 3206 7404
rect 4080 7392 4108 7432
rect 6454 7420 6460 7432
rect 6512 7420 6518 7472
rect 7374 7460 7380 7472
rect 6564 7432 7380 7460
rect 3200 7364 4108 7392
rect 4157 7395 4215 7401
rect 3200 7352 3206 7364
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4430 7392 4436 7404
rect 4387 7364 4436 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 3602 7284 3608 7336
rect 3660 7324 3666 7336
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 3660 7296 4077 7324
rect 3660 7284 3666 7296
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 4172 7324 4200 7355
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4798 7352 4804 7404
rect 4856 7352 4862 7404
rect 6564 7392 6592 7432
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 9324 7469 9352 7500
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 17034 7488 17040 7540
rect 17092 7528 17098 7540
rect 18322 7528 18328 7540
rect 17092 7500 18328 7528
rect 17092 7488 17098 7500
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 21542 7528 21548 7540
rect 18524 7500 21548 7528
rect 9309 7463 9367 7469
rect 9309 7429 9321 7463
rect 9355 7429 9367 7463
rect 9309 7423 9367 7429
rect 10410 7420 10416 7472
rect 10468 7460 10474 7472
rect 12069 7463 12127 7469
rect 12069 7460 12081 7463
rect 10468 7432 12081 7460
rect 10468 7420 10474 7432
rect 12069 7429 12081 7432
rect 12115 7429 12127 7463
rect 12069 7423 12127 7429
rect 12161 7463 12219 7469
rect 12161 7429 12173 7463
rect 12207 7460 12219 7463
rect 12710 7460 12716 7472
rect 12207 7432 12716 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 4908 7364 6592 7392
rect 4908 7324 4936 7364
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 10870 7392 10876 7404
rect 8510 7364 10876 7392
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7392 11023 7395
rect 11790 7392 11796 7404
rect 11011 7364 11796 7392
rect 11011 7361 11023 7364
rect 10965 7355 11023 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 4172 7296 4936 7324
rect 4065 7287 4123 7293
rect 5718 7284 5724 7336
rect 5776 7284 5782 7336
rect 5810 7284 5816 7336
rect 5868 7284 5874 7336
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 9122 7324 9128 7336
rect 7423 7296 9128 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 10045 7327 10103 7333
rect 10045 7324 10057 7327
rect 9364 7296 10057 7324
rect 9364 7284 9370 7296
rect 10045 7293 10057 7296
rect 10091 7293 10103 7327
rect 10045 7287 10103 7293
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 12176 7324 12204 7423
rect 12710 7420 12716 7432
rect 12768 7420 12774 7472
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 13081 7463 13139 7469
rect 13081 7460 13093 7463
rect 13044 7432 13093 7460
rect 13044 7420 13050 7432
rect 13081 7429 13093 7432
rect 13127 7429 13139 7463
rect 13081 7423 13139 7429
rect 14185 7463 14243 7469
rect 14185 7429 14197 7463
rect 14231 7460 14243 7463
rect 14458 7460 14464 7472
rect 14231 7432 14464 7460
rect 14231 7429 14243 7432
rect 14185 7423 14243 7429
rect 14458 7420 14464 7432
rect 14516 7420 14522 7472
rect 14734 7420 14740 7472
rect 14792 7420 14798 7472
rect 15933 7463 15991 7469
rect 15933 7429 15945 7463
rect 15979 7460 15991 7463
rect 16758 7460 16764 7472
rect 15979 7432 16764 7460
rect 15979 7429 15991 7432
rect 15933 7423 15991 7429
rect 16758 7420 16764 7432
rect 16816 7420 16822 7472
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 18524 7469 18552 7500
rect 21542 7488 21548 7500
rect 21600 7488 21606 7540
rect 23382 7488 23388 7540
rect 23440 7488 23446 7540
rect 23845 7531 23903 7537
rect 23845 7497 23857 7531
rect 23891 7528 23903 7531
rect 24118 7528 24124 7540
rect 23891 7500 24124 7528
rect 23891 7497 23903 7500
rect 23845 7491 23903 7497
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 24883 7531 24941 7537
rect 24883 7497 24895 7531
rect 24929 7528 24941 7531
rect 25682 7528 25688 7540
rect 24929 7500 25688 7528
rect 24929 7497 24941 7500
rect 24883 7491 24941 7497
rect 25682 7488 25688 7500
rect 25740 7528 25746 7540
rect 25866 7528 25872 7540
rect 25740 7500 25872 7528
rect 25740 7488 25746 7500
rect 25866 7488 25872 7500
rect 25924 7488 25930 7540
rect 26970 7488 26976 7540
rect 27028 7528 27034 7540
rect 27157 7531 27215 7537
rect 27157 7528 27169 7531
rect 27028 7500 27169 7528
rect 27028 7488 27034 7500
rect 27157 7497 27169 7500
rect 27203 7497 27215 7531
rect 27157 7491 27215 7497
rect 27338 7488 27344 7540
rect 27396 7528 27402 7540
rect 27617 7531 27675 7537
rect 27617 7528 27629 7531
rect 27396 7500 27629 7528
rect 27396 7488 27402 7500
rect 27617 7497 27629 7500
rect 27663 7497 27675 7531
rect 27617 7491 27675 7497
rect 28166 7488 28172 7540
rect 28224 7528 28230 7540
rect 30929 7531 30987 7537
rect 28224 7500 30604 7528
rect 28224 7488 28230 7500
rect 18509 7463 18567 7469
rect 18509 7460 18521 7463
rect 17000 7432 18521 7460
rect 17000 7420 17006 7432
rect 18509 7429 18521 7432
rect 18555 7429 18567 7463
rect 18725 7463 18783 7469
rect 18725 7460 18737 7463
rect 18509 7423 18567 7429
rect 18708 7429 18737 7460
rect 18771 7460 18783 7463
rect 18874 7460 18880 7472
rect 18771 7432 18880 7460
rect 18771 7429 18783 7432
rect 18708 7423 18783 7429
rect 12802 7352 12808 7404
rect 12860 7392 12866 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12860 7364 12909 7392
rect 12860 7352 12866 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13170 7352 13176 7404
rect 13228 7352 13234 7404
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 11296 7296 12204 7324
rect 12345 7327 12403 7333
rect 11296 7284 11302 7296
rect 12345 7293 12357 7327
rect 12391 7293 12403 7327
rect 12345 7287 12403 7293
rect 2774 7216 2780 7268
rect 2832 7256 2838 7268
rect 11057 7259 11115 7265
rect 2832 7228 7144 7256
rect 2832 7216 2838 7228
rect 5074 7188 5080 7200
rect 2700 7160 5080 7188
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 5258 7148 5264 7200
rect 5316 7148 5322 7200
rect 5626 7148 5632 7200
rect 5684 7188 5690 7200
rect 6270 7188 6276 7200
rect 5684 7160 6276 7188
rect 5684 7148 5690 7160
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 6822 7188 6828 7200
rect 6604 7160 6828 7188
rect 6604 7148 6610 7160
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 7116 7188 7144 7228
rect 11057 7225 11069 7259
rect 11103 7256 11115 7259
rect 12066 7256 12072 7268
rect 11103 7228 12072 7256
rect 11103 7225 11115 7228
rect 11057 7219 11115 7225
rect 12066 7216 12072 7228
rect 12124 7216 12130 7268
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 12360 7256 12388 7287
rect 12526 7284 12532 7336
rect 12584 7324 12590 7336
rect 13280 7324 13308 7355
rect 13722 7352 13728 7404
rect 13780 7392 13786 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13780 7364 13921 7392
rect 13780 7352 13786 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 17310 7352 17316 7404
rect 17368 7392 17374 7404
rect 17681 7395 17739 7401
rect 17681 7392 17693 7395
rect 17368 7364 17693 7392
rect 17368 7352 17374 7364
rect 17681 7361 17693 7364
rect 17727 7361 17739 7395
rect 17681 7355 17739 7361
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7392 17831 7395
rect 18598 7392 18604 7404
rect 17819 7364 18604 7392
rect 17819 7361 17831 7364
rect 17773 7355 17831 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 13446 7324 13452 7336
rect 12584 7296 13308 7324
rect 13372 7296 13452 7324
rect 12584 7284 12590 7296
rect 13372 7256 13400 7296
rect 13446 7284 13452 7296
rect 13504 7324 13510 7336
rect 17865 7327 17923 7333
rect 17865 7324 17877 7327
rect 13504 7296 17877 7324
rect 13504 7284 13510 7296
rect 17865 7293 17877 7296
rect 17911 7293 17923 7327
rect 17865 7287 17923 7293
rect 17954 7284 17960 7336
rect 18012 7324 18018 7336
rect 18708 7324 18736 7423
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 20990 7460 20996 7472
rect 20838 7432 20996 7460
rect 20990 7420 20996 7432
rect 21048 7420 21054 7472
rect 22462 7420 22468 7472
rect 22520 7460 22526 7472
rect 22557 7463 22615 7469
rect 22557 7460 22569 7463
rect 22520 7432 22569 7460
rect 22520 7420 22526 7432
rect 22557 7429 22569 7432
rect 22603 7460 22615 7463
rect 22603 7432 23244 7460
rect 22603 7429 22615 7432
rect 22557 7423 22615 7429
rect 19334 7352 19340 7404
rect 19392 7352 19398 7404
rect 22370 7352 22376 7404
rect 22428 7352 22434 7404
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 19613 7327 19671 7333
rect 19613 7324 19625 7327
rect 18012 7296 18736 7324
rect 19444 7296 19625 7324
rect 18012 7284 18018 7296
rect 17972 7256 18000 7284
rect 12308 7228 13400 7256
rect 15212 7228 18000 7256
rect 12308 7216 12314 7228
rect 8849 7191 8907 7197
rect 8849 7188 8861 7191
rect 7116 7160 8861 7188
rect 8849 7157 8861 7160
rect 8895 7188 8907 7191
rect 9582 7188 9588 7200
rect 8895 7160 9588 7188
rect 8895 7157 8907 7160
rect 8849 7151 8907 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 11698 7148 11704 7200
rect 11756 7148 11762 7200
rect 13449 7191 13507 7197
rect 13449 7157 13461 7191
rect 13495 7188 13507 7191
rect 13814 7188 13820 7200
rect 13495 7160 13820 7188
rect 13495 7157 13507 7160
rect 13449 7151 13507 7157
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 15212 7188 15240 7228
rect 18138 7216 18144 7268
rect 18196 7256 18202 7268
rect 19444 7256 19472 7296
rect 19613 7293 19625 7296
rect 19659 7293 19671 7327
rect 19613 7287 19671 7293
rect 20806 7284 20812 7336
rect 20864 7324 20870 7336
rect 21361 7327 21419 7333
rect 21361 7324 21373 7327
rect 20864 7296 21373 7324
rect 20864 7284 20870 7296
rect 21361 7293 21373 7296
rect 21407 7293 21419 7327
rect 21361 7287 21419 7293
rect 21450 7284 21456 7336
rect 21508 7324 21514 7336
rect 22664 7324 22692 7355
rect 22738 7352 22744 7404
rect 22796 7352 22802 7404
rect 23216 7392 23244 7432
rect 23290 7420 23296 7472
rect 23348 7460 23354 7472
rect 24673 7463 24731 7469
rect 24673 7460 24685 7463
rect 23348 7432 24685 7460
rect 23348 7420 23354 7432
rect 24673 7429 24685 7432
rect 24719 7429 24731 7463
rect 25222 7460 25228 7472
rect 24673 7423 24731 7429
rect 24964 7432 25228 7460
rect 23216 7364 23704 7392
rect 21508 7296 22692 7324
rect 21508 7284 21514 7296
rect 18196 7228 19472 7256
rect 23676 7256 23704 7364
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 24486 7392 24492 7404
rect 23808 7364 24492 7392
rect 23808 7352 23814 7364
rect 24486 7352 24492 7364
rect 24544 7352 24550 7404
rect 24964 7392 24992 7432
rect 25222 7420 25228 7432
rect 25280 7420 25286 7472
rect 25498 7420 25504 7472
rect 25556 7420 25562 7472
rect 27525 7463 27583 7469
rect 27525 7429 27537 7463
rect 27571 7460 27583 7463
rect 27982 7460 27988 7472
rect 27571 7432 27988 7460
rect 27571 7429 27583 7432
rect 27525 7423 27583 7429
rect 27982 7420 27988 7432
rect 28040 7420 28046 7472
rect 28994 7460 29000 7472
rect 28644 7432 29000 7460
rect 24964 7364 25084 7392
rect 24029 7327 24087 7333
rect 24029 7293 24041 7327
rect 24075 7324 24087 7327
rect 24854 7324 24860 7336
rect 24075 7296 24860 7324
rect 24075 7293 24087 7296
rect 24029 7287 24087 7293
rect 24854 7284 24860 7296
rect 24912 7284 24918 7336
rect 25056 7265 25084 7364
rect 25958 7352 25964 7404
rect 26016 7392 26022 7404
rect 28350 7392 28356 7404
rect 26016 7364 28356 7392
rect 26016 7352 26022 7364
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 28644 7401 28672 7432
rect 28994 7420 29000 7432
rect 29052 7420 29058 7472
rect 29362 7420 29368 7472
rect 29420 7420 29426 7472
rect 28629 7395 28687 7401
rect 28629 7361 28641 7395
rect 28675 7361 28687 7395
rect 30576 7392 30604 7500
rect 30929 7497 30941 7531
rect 30975 7528 30987 7531
rect 31018 7528 31024 7540
rect 30975 7500 31024 7528
rect 30975 7497 30987 7500
rect 30929 7491 30987 7497
rect 31018 7488 31024 7500
rect 31076 7488 31082 7540
rect 31297 7531 31355 7537
rect 31297 7497 31309 7531
rect 31343 7528 31355 7531
rect 32398 7528 32404 7540
rect 31343 7500 32404 7528
rect 31343 7497 31355 7500
rect 31297 7491 31355 7497
rect 31312 7460 31340 7491
rect 32398 7488 32404 7500
rect 32456 7488 32462 7540
rect 32674 7488 32680 7540
rect 32732 7528 32738 7540
rect 34267 7531 34325 7537
rect 34267 7528 34279 7531
rect 32732 7500 34279 7528
rect 32732 7488 32738 7500
rect 34267 7497 34279 7500
rect 34313 7528 34325 7531
rect 35250 7528 35256 7540
rect 34313 7500 35256 7528
rect 34313 7497 34325 7500
rect 34267 7491 34325 7497
rect 35250 7488 35256 7500
rect 35308 7488 35314 7540
rect 36170 7528 36176 7540
rect 35360 7500 36176 7528
rect 30839 7432 31340 7460
rect 30839 7392 30867 7432
rect 34054 7420 34060 7472
rect 34112 7420 34118 7472
rect 35360 7460 35388 7500
rect 36170 7488 36176 7500
rect 36228 7488 36234 7540
rect 36906 7488 36912 7540
rect 36964 7488 36970 7540
rect 37182 7488 37188 7540
rect 37240 7528 37246 7540
rect 37829 7531 37887 7537
rect 37829 7528 37841 7531
rect 37240 7500 37841 7528
rect 37240 7488 37246 7500
rect 37829 7497 37841 7500
rect 37875 7497 37887 7531
rect 37829 7491 37887 7497
rect 35176 7432 35388 7460
rect 30576 7364 30867 7392
rect 31389 7395 31447 7401
rect 28629 7355 28687 7361
rect 31389 7361 31401 7395
rect 31435 7392 31447 7395
rect 31754 7392 31760 7404
rect 31435 7364 31760 7392
rect 31435 7361 31447 7364
rect 31389 7355 31447 7361
rect 31754 7352 31760 7364
rect 31812 7352 31818 7404
rect 32674 7352 32680 7404
rect 32732 7352 32738 7404
rect 33226 7352 33232 7404
rect 33284 7392 33290 7404
rect 35176 7401 35204 7432
rect 35986 7420 35992 7472
rect 36044 7420 36050 7472
rect 36924 7460 36952 7488
rect 37921 7463 37979 7469
rect 37921 7460 37933 7463
rect 36924 7432 37933 7460
rect 37921 7429 37933 7432
rect 37967 7429 37979 7463
rect 37921 7423 37979 7429
rect 33505 7395 33563 7401
rect 33505 7392 33517 7395
rect 33284 7364 33517 7392
rect 33284 7352 33290 7364
rect 33505 7361 33517 7364
rect 33551 7392 33563 7395
rect 35161 7395 35219 7401
rect 35161 7392 35173 7395
rect 33551 7364 35173 7392
rect 33551 7361 33563 7364
rect 33505 7355 33563 7361
rect 35161 7361 35173 7364
rect 35207 7361 35219 7395
rect 35161 7355 35219 7361
rect 25130 7284 25136 7336
rect 25188 7324 25194 7336
rect 26237 7327 26295 7333
rect 26237 7324 26249 7327
rect 25188 7296 26249 7324
rect 25188 7284 25194 7296
rect 26237 7293 26249 7296
rect 26283 7324 26295 7327
rect 26786 7324 26792 7336
rect 26283 7296 26792 7324
rect 26283 7293 26295 7296
rect 26237 7287 26295 7293
rect 26786 7284 26792 7296
rect 26844 7284 26850 7336
rect 27709 7327 27767 7333
rect 27709 7293 27721 7327
rect 27755 7293 27767 7327
rect 27709 7287 27767 7293
rect 25041 7259 25099 7265
rect 23676 7228 24992 7256
rect 18196 7216 18202 7228
rect 14332 7160 15240 7188
rect 14332 7148 14338 7160
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 17126 7188 17132 7200
rect 16448 7160 17132 7188
rect 16448 7148 16454 7160
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 17313 7191 17371 7197
rect 17313 7157 17325 7191
rect 17359 7188 17371 7191
rect 17402 7188 17408 7200
rect 17359 7160 17408 7188
rect 17359 7157 17371 7160
rect 17313 7151 17371 7157
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 18693 7191 18751 7197
rect 18693 7188 18705 7191
rect 17920 7160 18705 7188
rect 17920 7148 17926 7160
rect 18693 7157 18705 7160
rect 18739 7157 18751 7191
rect 18693 7151 18751 7157
rect 18877 7191 18935 7197
rect 18877 7157 18889 7191
rect 18923 7188 18935 7191
rect 21082 7188 21088 7200
rect 18923 7160 21088 7188
rect 18923 7157 18935 7160
rect 18877 7151 18935 7157
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 21174 7148 21180 7200
rect 21232 7188 21238 7200
rect 22925 7191 22983 7197
rect 22925 7188 22937 7191
rect 21232 7160 22937 7188
rect 21232 7148 21238 7160
rect 22925 7157 22937 7160
rect 22971 7157 22983 7191
rect 22925 7151 22983 7157
rect 24854 7148 24860 7200
rect 24912 7148 24918 7200
rect 24964 7188 24992 7228
rect 25041 7225 25053 7259
rect 25087 7225 25099 7259
rect 25041 7219 25099 7225
rect 25774 7216 25780 7268
rect 25832 7256 25838 7268
rect 27724 7256 27752 7287
rect 27798 7284 27804 7336
rect 27856 7324 27862 7336
rect 28905 7327 28963 7333
rect 28905 7324 28917 7327
rect 27856 7296 28917 7324
rect 27856 7284 27862 7296
rect 28905 7293 28917 7296
rect 28951 7293 28963 7327
rect 28905 7287 28963 7293
rect 30282 7284 30288 7336
rect 30340 7324 30346 7336
rect 30377 7327 30435 7333
rect 30377 7324 30389 7327
rect 30340 7296 30389 7324
rect 30340 7284 30346 7296
rect 30377 7293 30389 7296
rect 30423 7293 30435 7327
rect 30377 7287 30435 7293
rect 31202 7284 31208 7336
rect 31260 7324 31266 7336
rect 31570 7324 31576 7336
rect 31260 7296 31576 7324
rect 31260 7284 31266 7296
rect 31570 7284 31576 7296
rect 31628 7284 31634 7336
rect 32398 7284 32404 7336
rect 32456 7324 32462 7336
rect 34698 7324 34704 7336
rect 32456 7296 34704 7324
rect 32456 7284 32462 7296
rect 34698 7284 34704 7296
rect 34756 7284 34762 7336
rect 35437 7327 35495 7333
rect 35437 7293 35449 7327
rect 35483 7324 35495 7327
rect 35483 7296 37504 7324
rect 35483 7293 35495 7296
rect 35437 7287 35495 7293
rect 31386 7256 31392 7268
rect 25832 7228 27752 7256
rect 25832 7216 25838 7228
rect 25958 7188 25964 7200
rect 24964 7160 25964 7188
rect 25958 7148 25964 7160
rect 26016 7148 26022 7200
rect 27724 7188 27752 7228
rect 30208 7228 31392 7256
rect 30208 7188 30236 7228
rect 31386 7216 31392 7228
rect 31444 7216 31450 7268
rect 37476 7265 37504 7296
rect 37734 7284 37740 7336
rect 37792 7324 37798 7336
rect 38013 7327 38071 7333
rect 38013 7324 38025 7327
rect 37792 7296 38025 7324
rect 37792 7284 37798 7296
rect 38013 7293 38025 7296
rect 38059 7293 38071 7327
rect 38013 7287 38071 7293
rect 34425 7259 34483 7265
rect 34425 7256 34437 7259
rect 31588 7228 34437 7256
rect 27724 7160 30236 7188
rect 30282 7148 30288 7200
rect 30340 7188 30346 7200
rect 31588 7188 31616 7228
rect 34425 7225 34437 7228
rect 34471 7225 34483 7259
rect 34425 7219 34483 7225
rect 37461 7259 37519 7265
rect 37461 7225 37473 7259
rect 37507 7225 37519 7259
rect 37461 7219 37519 7225
rect 30340 7160 31616 7188
rect 30340 7148 30346 7160
rect 31662 7148 31668 7200
rect 31720 7188 31726 7200
rect 34241 7191 34299 7197
rect 34241 7188 34253 7191
rect 31720 7160 34253 7188
rect 31720 7148 31726 7160
rect 34241 7157 34253 7160
rect 34287 7188 34299 7191
rect 36722 7188 36728 7200
rect 34287 7160 36728 7188
rect 34287 7157 34299 7160
rect 34241 7151 34299 7157
rect 36722 7148 36728 7160
rect 36780 7148 36786 7200
rect 1104 7098 39192 7120
rect 1104 7046 5711 7098
rect 5763 7046 5775 7098
rect 5827 7046 5839 7098
rect 5891 7046 5903 7098
rect 5955 7046 5967 7098
rect 6019 7046 15233 7098
rect 15285 7046 15297 7098
rect 15349 7046 15361 7098
rect 15413 7046 15425 7098
rect 15477 7046 15489 7098
rect 15541 7046 24755 7098
rect 24807 7046 24819 7098
rect 24871 7046 24883 7098
rect 24935 7046 24947 7098
rect 24999 7046 25011 7098
rect 25063 7046 34277 7098
rect 34329 7046 34341 7098
rect 34393 7046 34405 7098
rect 34457 7046 34469 7098
rect 34521 7046 34533 7098
rect 34585 7046 39192 7098
rect 1104 7024 39192 7046
rect 2041 6987 2099 6993
rect 2041 6953 2053 6987
rect 2087 6984 2099 6987
rect 2958 6984 2964 6996
rect 2087 6956 2964 6984
rect 2087 6953 2099 6956
rect 2041 6947 2099 6953
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 5432 6987 5490 6993
rect 5432 6953 5444 6987
rect 5478 6984 5490 6987
rect 11698 6984 11704 6996
rect 5478 6956 11704 6984
rect 5478 6953 5490 6956
rect 5432 6947 5490 6953
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 14734 6984 14740 6996
rect 12124 6956 14740 6984
rect 12124 6944 12130 6956
rect 14734 6944 14740 6956
rect 14792 6944 14798 6996
rect 15102 6944 15108 6996
rect 15160 6984 15166 6996
rect 15160 6956 15884 6984
rect 15160 6944 15166 6956
rect 4430 6876 4436 6928
rect 4488 6916 4494 6928
rect 12805 6919 12863 6925
rect 4488 6888 4660 6916
rect 4488 6876 4494 6888
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 3329 6851 3387 6857
rect 1912 6820 2774 6848
rect 1912 6808 1918 6820
rect 2746 6780 2774 6820
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 4338 6848 4344 6860
rect 3375 6820 4344 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 4632 6857 4660 6888
rect 12805 6885 12817 6919
rect 12851 6916 12863 6919
rect 12894 6916 12900 6928
rect 12851 6888 12900 6916
rect 12851 6885 12863 6888
rect 12805 6879 12863 6885
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 13630 6876 13636 6928
rect 13688 6916 13694 6928
rect 14274 6916 14280 6928
rect 13688 6888 14280 6916
rect 13688 6876 13694 6888
rect 14274 6876 14280 6888
rect 14332 6876 14338 6928
rect 15378 6876 15384 6928
rect 15436 6916 15442 6928
rect 15746 6916 15752 6928
rect 15436 6888 15752 6916
rect 15436 6876 15442 6888
rect 15746 6876 15752 6888
rect 15804 6876 15810 6928
rect 15856 6916 15884 6956
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 17018 6987 17076 6993
rect 17018 6984 17030 6987
rect 15988 6956 17030 6984
rect 15988 6944 15994 6956
rect 17018 6953 17030 6956
rect 17064 6953 17076 6987
rect 17018 6947 17076 6953
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17184 6956 18092 6984
rect 17184 6944 17190 6956
rect 16666 6916 16672 6928
rect 15856 6888 16672 6916
rect 16666 6876 16672 6888
rect 16724 6916 16730 6928
rect 18064 6916 18092 6956
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 20806 6984 20812 6996
rect 18380 6956 20812 6984
rect 18380 6944 18386 6956
rect 20806 6944 20812 6956
rect 20864 6944 20870 6996
rect 21082 6944 21088 6996
rect 21140 6944 21146 6996
rect 22268 6987 22326 6993
rect 22268 6953 22280 6987
rect 22314 6984 22326 6987
rect 25222 6984 25228 6996
rect 22314 6956 25228 6984
rect 22314 6953 22326 6956
rect 22268 6947 22326 6953
rect 25222 6944 25228 6956
rect 25280 6944 25286 6996
rect 26142 6944 26148 6996
rect 26200 6984 26206 6996
rect 26970 6984 26976 6996
rect 26200 6956 26976 6984
rect 26200 6944 26206 6956
rect 26970 6944 26976 6956
rect 27028 6944 27034 6996
rect 27154 6944 27160 6996
rect 27212 6984 27218 6996
rect 28721 6987 28779 6993
rect 28721 6984 28733 6987
rect 27212 6956 28733 6984
rect 27212 6944 27218 6956
rect 28721 6953 28733 6956
rect 28767 6953 28779 6987
rect 28721 6947 28779 6953
rect 28994 6944 29000 6996
rect 29052 6984 29058 6996
rect 31662 6984 31668 6996
rect 29052 6956 31668 6984
rect 29052 6944 29058 6956
rect 31662 6944 31668 6956
rect 31720 6944 31726 6996
rect 34149 6987 34207 6993
rect 34149 6953 34161 6987
rect 34195 6984 34207 6987
rect 35986 6984 35992 6996
rect 34195 6956 35992 6984
rect 34195 6953 34207 6956
rect 34149 6947 34207 6953
rect 35986 6944 35992 6956
rect 36044 6944 36050 6996
rect 36078 6944 36084 6996
rect 36136 6984 36142 6996
rect 37074 6987 37132 6993
rect 37074 6984 37086 6987
rect 36136 6956 37086 6984
rect 36136 6944 36142 6956
rect 37074 6953 37086 6956
rect 37120 6953 37132 6987
rect 37074 6947 37132 6953
rect 16724 6888 16804 6916
rect 18064 6888 18828 6916
rect 16724 6876 16730 6888
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 4798 6848 4804 6860
rect 4663 6820 4804 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6848 5227 6851
rect 6454 6848 6460 6860
rect 5215 6820 6460 6848
rect 5215 6817 5227 6820
rect 5169 6811 5227 6817
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 10502 6808 10508 6860
rect 10560 6808 10566 6860
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 11020 6820 11069 6848
rect 11020 6808 11026 6820
rect 11057 6817 11069 6820
rect 11103 6848 11115 6851
rect 13722 6848 13728 6860
rect 11103 6820 13728 6848
rect 11103 6817 11115 6820
rect 11057 6811 11115 6817
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 14369 6851 14427 6857
rect 14369 6817 14381 6851
rect 14415 6848 14427 6851
rect 16390 6848 16396 6860
rect 14415 6820 16396 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 16776 6857 16804 6888
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6817 16819 6851
rect 16761 6811 16819 6817
rect 18230 6808 18236 6860
rect 18288 6848 18294 6860
rect 18690 6848 18696 6860
rect 18288 6820 18696 6848
rect 18288 6808 18294 6820
rect 18690 6808 18696 6820
rect 18748 6808 18754 6860
rect 18800 6848 18828 6888
rect 19334 6876 19340 6928
rect 19392 6916 19398 6928
rect 19392 6888 22048 6916
rect 19392 6876 19398 6888
rect 20438 6848 20444 6860
rect 18800 6820 20444 6848
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 22020 6857 22048 6888
rect 26602 6876 26608 6928
rect 26660 6916 26666 6928
rect 26660 6888 28120 6916
rect 26660 6876 26666 6888
rect 22005 6851 22063 6857
rect 22005 6817 22017 6851
rect 22051 6848 22063 6851
rect 23658 6848 23664 6860
rect 22051 6820 23664 6848
rect 22051 6817 22063 6820
rect 22005 6811 22063 6817
rect 23658 6808 23664 6820
rect 23716 6848 23722 6860
rect 25130 6848 25136 6860
rect 23716 6820 25136 6848
rect 23716 6808 23722 6820
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 25406 6808 25412 6860
rect 25464 6848 25470 6860
rect 27157 6851 27215 6857
rect 27157 6848 27169 6851
rect 25464 6820 27169 6848
rect 25464 6808 25470 6820
rect 27157 6817 27169 6820
rect 27203 6817 27215 6851
rect 27157 6811 27215 6817
rect 4430 6780 4436 6792
rect 2746 6752 4436 6780
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 7650 6740 7656 6792
rect 7708 6740 7714 6792
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 9766 6780 9772 6792
rect 9263 6752 9772 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 10192 6752 10241 6780
rect 10192 6740 10198 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 13044 6752 13277 6780
rect 13044 6740 13050 6752
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 14056 6752 14289 6780
rect 14056 6740 14062 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14921 6783 14979 6789
rect 14921 6749 14933 6783
rect 14967 6780 14979 6783
rect 15010 6780 15016 6792
rect 14967 6752 15016 6780
rect 14967 6749 14979 6752
rect 14921 6743 14979 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 20257 6783 20315 6789
rect 20257 6780 20269 6783
rect 19576 6752 20269 6780
rect 19576 6740 19582 6752
rect 20257 6749 20269 6752
rect 20303 6780 20315 6783
rect 20530 6780 20536 6792
rect 20303 6752 20536 6780
rect 20303 6749 20315 6752
rect 20257 6743 20315 6749
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 21082 6740 21088 6792
rect 21140 6740 21146 6792
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 27522 6780 27528 6792
rect 26542 6752 27528 6780
rect 21177 6743 21235 6749
rect 1857 6715 1915 6721
rect 1857 6681 1869 6715
rect 1903 6712 1915 6715
rect 1946 6712 1952 6724
rect 1903 6684 1952 6712
rect 1903 6681 1915 6684
rect 1857 6675 1915 6681
rect 1946 6672 1952 6684
rect 2004 6672 2010 6724
rect 2130 6721 2136 6724
rect 2073 6715 2136 6721
rect 2073 6681 2085 6715
rect 2119 6681 2136 6715
rect 2073 6675 2136 6681
rect 2130 6672 2136 6675
rect 2188 6672 2194 6724
rect 2406 6712 2412 6724
rect 2240 6684 2412 6712
rect 2240 6653 2268 6684
rect 2406 6672 2412 6684
rect 2464 6672 2470 6724
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 2866 6712 2872 6724
rect 2648 6684 2872 6712
rect 2648 6672 2654 6684
rect 2866 6672 2872 6684
rect 2924 6672 2930 6724
rect 3053 6715 3111 6721
rect 3053 6681 3065 6715
rect 3099 6712 3111 6715
rect 4154 6712 4160 6724
rect 3099 6684 4160 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 4304 6684 4476 6712
rect 4304 6672 4310 6684
rect 2225 6647 2283 6653
rect 2225 6613 2237 6647
rect 2271 6613 2283 6647
rect 2225 6607 2283 6613
rect 2314 6604 2320 6656
rect 2372 6644 2378 6656
rect 2685 6647 2743 6653
rect 2685 6644 2697 6647
rect 2372 6616 2697 6644
rect 2372 6604 2378 6616
rect 2685 6613 2697 6616
rect 2731 6613 2743 6647
rect 2685 6607 2743 6613
rect 3142 6604 3148 6656
rect 3200 6604 3206 6656
rect 3970 6604 3976 6656
rect 4028 6604 4034 6656
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4448 6653 4476 6684
rect 6454 6672 6460 6724
rect 6512 6672 6518 6724
rect 7006 6712 7012 6724
rect 6748 6684 7012 6712
rect 4341 6647 4399 6653
rect 4341 6644 4353 6647
rect 4120 6616 4353 6644
rect 4120 6604 4126 6616
rect 4341 6613 4353 6616
rect 4387 6613 4399 6647
rect 4341 6607 4399 6613
rect 4433 6647 4491 6653
rect 4433 6613 4445 6647
rect 4479 6613 4491 6647
rect 4433 6607 4491 6613
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6748 6644 6776 6684
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 8386 6672 8392 6724
rect 8444 6672 8450 6724
rect 11238 6712 11244 6724
rect 9232 6684 11244 6712
rect 5592 6616 6776 6644
rect 6917 6647 6975 6653
rect 5592 6604 5598 6616
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 9232 6644 9260 6684
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 11330 6672 11336 6724
rect 11388 6672 11394 6724
rect 13541 6715 13599 6721
rect 12728 6684 13492 6712
rect 6963 6616 9260 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 9306 6604 9312 6656
rect 9364 6604 9370 6656
rect 9858 6604 9864 6656
rect 9916 6604 9922 6656
rect 10321 6647 10379 6653
rect 10321 6613 10333 6647
rect 10367 6644 10379 6647
rect 12728 6644 12756 6684
rect 10367 6616 12756 6644
rect 13464 6644 13492 6684
rect 13541 6681 13553 6715
rect 13587 6712 13599 6715
rect 15378 6712 15384 6724
rect 13587 6684 15384 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 15378 6672 15384 6684
rect 15436 6672 15442 6724
rect 15470 6672 15476 6724
rect 15528 6712 15534 6724
rect 15657 6715 15715 6721
rect 15657 6712 15669 6715
rect 15528 6684 15669 6712
rect 15528 6672 15534 6684
rect 15657 6681 15669 6684
rect 15703 6681 15715 6715
rect 16942 6712 16948 6724
rect 15657 6675 15715 6681
rect 15856 6684 16948 6712
rect 15856 6644 15884 6684
rect 16942 6672 16948 6684
rect 17000 6672 17006 6724
rect 17494 6672 17500 6724
rect 17552 6672 17558 6724
rect 18782 6672 18788 6724
rect 18840 6672 18846 6724
rect 19702 6672 19708 6724
rect 19760 6712 19766 6724
rect 20349 6715 20407 6721
rect 20349 6712 20361 6715
rect 19760 6684 20361 6712
rect 19760 6672 19766 6684
rect 20349 6681 20361 6684
rect 20395 6681 20407 6715
rect 20349 6675 20407 6681
rect 20622 6672 20628 6724
rect 20680 6712 20686 6724
rect 21192 6712 21220 6743
rect 27522 6740 27528 6752
rect 27580 6740 27586 6792
rect 27614 6740 27620 6792
rect 27672 6740 27678 6792
rect 27798 6789 27804 6792
rect 27765 6783 27804 6789
rect 27765 6749 27777 6783
rect 27765 6743 27804 6749
rect 27798 6740 27804 6743
rect 27856 6740 27862 6792
rect 27982 6740 27988 6792
rect 28040 6740 28046 6792
rect 28092 6789 28120 6888
rect 28258 6876 28264 6928
rect 28316 6916 28322 6928
rect 31386 6916 31392 6928
rect 28316 6888 31392 6916
rect 28316 6876 28322 6888
rect 31386 6876 31392 6888
rect 31444 6876 31450 6928
rect 31478 6876 31484 6928
rect 31536 6916 31542 6928
rect 34882 6916 34888 6928
rect 31536 6888 34888 6916
rect 31536 6876 31542 6888
rect 34882 6876 34888 6888
rect 34940 6916 34946 6928
rect 34940 6888 35480 6916
rect 34940 6876 34946 6888
rect 28905 6851 28963 6857
rect 28905 6817 28917 6851
rect 28951 6848 28963 6851
rect 30282 6848 30288 6860
rect 28951 6820 30288 6848
rect 28951 6817 28963 6820
rect 28905 6811 28963 6817
rect 30282 6808 30288 6820
rect 30340 6808 30346 6860
rect 30742 6808 30748 6860
rect 30800 6848 30806 6860
rect 30929 6851 30987 6857
rect 30929 6848 30941 6851
rect 30800 6820 30941 6848
rect 30800 6808 30806 6820
rect 30929 6817 30941 6820
rect 30975 6817 30987 6851
rect 30929 6811 30987 6817
rect 31113 6851 31171 6857
rect 31113 6817 31125 6851
rect 31159 6817 31171 6851
rect 31113 6811 31171 6817
rect 28082 6783 28140 6789
rect 28082 6749 28094 6783
rect 28128 6749 28140 6783
rect 28082 6743 28140 6749
rect 28258 6740 28264 6792
rect 28316 6740 28322 6792
rect 28997 6783 29055 6789
rect 28997 6749 29009 6783
rect 29043 6780 29055 6783
rect 29270 6780 29276 6792
rect 29043 6752 29276 6780
rect 29043 6749 29055 6752
rect 28997 6743 29055 6749
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 31128 6780 31156 6811
rect 31294 6808 31300 6860
rect 31352 6848 31358 6860
rect 35452 6857 35480 6888
rect 35437 6851 35495 6857
rect 31352 6820 32812 6848
rect 31352 6808 31358 6820
rect 31478 6780 31484 6792
rect 29748 6752 31064 6780
rect 31128 6752 31484 6780
rect 20680 6684 21220 6712
rect 20680 6672 20686 6684
rect 22922 6672 22928 6724
rect 22980 6672 22986 6724
rect 24029 6715 24087 6721
rect 24029 6681 24041 6715
rect 24075 6681 24087 6715
rect 24029 6675 24087 6681
rect 13464 6616 15884 6644
rect 10367 6613 10379 6616
rect 10321 6607 10379 6613
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 19889 6647 19947 6653
rect 19889 6644 19901 6647
rect 15988 6616 19901 6644
rect 15988 6604 15994 6616
rect 19889 6613 19901 6616
rect 19935 6613 19947 6647
rect 19889 6607 19947 6613
rect 21450 6604 21456 6656
rect 21508 6604 21514 6656
rect 24044 6644 24072 6675
rect 25406 6672 25412 6724
rect 25464 6672 25470 6724
rect 27338 6672 27344 6724
rect 27396 6712 27402 6724
rect 27893 6715 27951 6721
rect 27893 6712 27905 6715
rect 27396 6684 27905 6712
rect 27396 6672 27402 6684
rect 27893 6681 27905 6684
rect 27939 6712 27951 6715
rect 28276 6712 28304 6740
rect 27939 6684 28304 6712
rect 28721 6715 28779 6721
rect 27939 6681 27951 6684
rect 27893 6675 27951 6681
rect 28721 6681 28733 6715
rect 28767 6712 28779 6715
rect 29748 6712 29776 6752
rect 28767 6684 29776 6712
rect 29825 6715 29883 6721
rect 28767 6681 28779 6684
rect 28721 6675 28779 6681
rect 29825 6681 29837 6715
rect 29871 6681 29883 6715
rect 29825 6675 29883 6681
rect 30837 6715 30895 6721
rect 30837 6681 30849 6715
rect 30883 6712 30895 6715
rect 30926 6712 30932 6724
rect 30883 6684 30932 6712
rect 30883 6681 30895 6684
rect 30837 6675 30895 6681
rect 28166 6644 28172 6656
rect 24044 6616 28172 6644
rect 28166 6604 28172 6616
rect 28224 6604 28230 6656
rect 28258 6604 28264 6656
rect 28316 6604 28322 6656
rect 29181 6647 29239 6653
rect 29181 6613 29193 6647
rect 29227 6644 29239 6647
rect 29840 6644 29868 6675
rect 30926 6672 30932 6684
rect 30984 6672 30990 6724
rect 29227 6616 29868 6644
rect 29227 6613 29239 6616
rect 29181 6607 29239 6613
rect 29914 6604 29920 6656
rect 29972 6604 29978 6656
rect 30466 6604 30472 6656
rect 30524 6604 30530 6656
rect 31036 6644 31064 6752
rect 31478 6740 31484 6752
rect 31536 6740 31542 6792
rect 31662 6740 31668 6792
rect 31720 6740 31726 6792
rect 31846 6740 31852 6792
rect 31904 6740 31910 6792
rect 32030 6740 32036 6792
rect 32088 6740 32094 6792
rect 32674 6740 32680 6792
rect 32732 6740 32738 6792
rect 32784 6780 32812 6820
rect 35437 6817 35449 6851
rect 35483 6848 35495 6851
rect 37734 6848 37740 6860
rect 35483 6820 37740 6848
rect 35483 6817 35495 6820
rect 35437 6811 35495 6817
rect 37734 6808 37740 6820
rect 37792 6808 37798 6860
rect 32784 6752 33640 6780
rect 31941 6715 31999 6721
rect 31941 6681 31953 6715
rect 31987 6712 31999 6715
rect 32766 6712 32772 6724
rect 31987 6684 32772 6712
rect 31987 6681 31999 6684
rect 31941 6675 31999 6681
rect 32766 6672 32772 6684
rect 32824 6672 32830 6724
rect 33502 6672 33508 6724
rect 33560 6672 33566 6724
rect 33612 6712 33640 6752
rect 34054 6740 34060 6792
rect 34112 6740 34118 6792
rect 34698 6740 34704 6792
rect 34756 6780 34762 6792
rect 35345 6783 35403 6789
rect 35345 6780 35357 6783
rect 34756 6752 35357 6780
rect 34756 6740 34762 6752
rect 35345 6749 35357 6752
rect 35391 6749 35403 6783
rect 35345 6743 35403 6749
rect 35802 6740 35808 6792
rect 35860 6780 35866 6792
rect 35986 6780 35992 6792
rect 35860 6752 35992 6780
rect 35860 6740 35866 6752
rect 35986 6740 35992 6752
rect 36044 6740 36050 6792
rect 36078 6740 36084 6792
rect 36136 6740 36142 6792
rect 36814 6740 36820 6792
rect 36872 6740 36878 6792
rect 36173 6715 36231 6721
rect 36173 6712 36185 6715
rect 33612 6684 34100 6712
rect 32217 6647 32275 6653
rect 32217 6644 32229 6647
rect 31036 6616 32229 6644
rect 32217 6613 32229 6616
rect 32263 6613 32275 6647
rect 34072 6644 34100 6684
rect 34256 6684 36185 6712
rect 34256 6644 34284 6684
rect 36173 6681 36185 6684
rect 36219 6681 36231 6715
rect 36173 6675 36231 6681
rect 37366 6672 37372 6724
rect 37424 6712 37430 6724
rect 37424 6684 37582 6712
rect 37424 6672 37430 6684
rect 34072 6616 34284 6644
rect 32217 6607 32275 6613
rect 34882 6604 34888 6656
rect 34940 6604 34946 6656
rect 35250 6604 35256 6656
rect 35308 6644 35314 6656
rect 37826 6644 37832 6656
rect 35308 6616 37832 6644
rect 35308 6604 35314 6616
rect 37826 6604 37832 6616
rect 37884 6604 37890 6656
rect 38562 6604 38568 6656
rect 38620 6604 38626 6656
rect 1104 6554 39352 6576
rect 1104 6502 10472 6554
rect 10524 6502 10536 6554
rect 10588 6502 10600 6554
rect 10652 6502 10664 6554
rect 10716 6502 10728 6554
rect 10780 6502 19994 6554
rect 20046 6502 20058 6554
rect 20110 6502 20122 6554
rect 20174 6502 20186 6554
rect 20238 6502 20250 6554
rect 20302 6502 29516 6554
rect 29568 6502 29580 6554
rect 29632 6502 29644 6554
rect 29696 6502 29708 6554
rect 29760 6502 29772 6554
rect 29824 6502 39038 6554
rect 39090 6502 39102 6554
rect 39154 6502 39166 6554
rect 39218 6502 39230 6554
rect 39282 6502 39294 6554
rect 39346 6502 39352 6554
rect 1104 6480 39352 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 3418 6440 3424 6452
rect 1811 6412 3424 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 4304 6412 5457 6440
rect 4304 6400 4310 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 6564 6412 6776 6440
rect 2685 6375 2743 6381
rect 2685 6341 2697 6375
rect 2731 6372 2743 6375
rect 3326 6372 3332 6384
rect 2731 6344 3332 6372
rect 2731 6341 2743 6344
rect 2685 6335 2743 6341
rect 3326 6332 3332 6344
rect 3384 6332 3390 6384
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 4430 6332 4436 6384
rect 4488 6332 4494 6384
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 6564 6372 6592 6412
rect 6748 6381 6776 6412
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7101 6443 7159 6449
rect 7101 6440 7113 6443
rect 6972 6412 7113 6440
rect 6972 6400 6978 6412
rect 7101 6409 7113 6412
rect 7147 6409 7159 6443
rect 7101 6403 7159 6409
rect 8018 6400 8024 6452
rect 8076 6400 8082 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10778 6440 10784 6452
rect 10284 6412 10784 6440
rect 10284 6400 10290 6412
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 12526 6400 12532 6452
rect 12584 6400 12590 6452
rect 12621 6443 12679 6449
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 13538 6440 13544 6452
rect 12667 6412 13544 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 6512 6344 6592 6372
rect 6733 6375 6791 6381
rect 6512 6332 6518 6344
rect 6733 6341 6745 6375
rect 6779 6372 6791 6375
rect 8036 6372 8064 6400
rect 6779 6344 8064 6372
rect 6779 6341 6791 6344
rect 6733 6335 6791 6341
rect 8294 6332 8300 6384
rect 8352 6332 8358 6384
rect 9585 6375 9643 6381
rect 9585 6341 9597 6375
rect 9631 6372 9643 6375
rect 12636 6372 12664 6403
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 13725 6443 13783 6449
rect 13725 6409 13737 6443
rect 13771 6440 13783 6443
rect 17218 6440 17224 6452
rect 13771 6412 17224 6440
rect 13771 6409 13783 6412
rect 13725 6403 13783 6409
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 22554 6440 22560 6452
rect 18012 6412 22560 6440
rect 18012 6400 18018 6412
rect 22554 6400 22560 6412
rect 22612 6400 22618 6452
rect 22830 6400 22836 6452
rect 22888 6440 22894 6452
rect 23385 6443 23443 6449
rect 23385 6440 23397 6443
rect 22888 6412 23397 6440
rect 22888 6400 22894 6412
rect 23385 6409 23397 6412
rect 23431 6409 23443 6443
rect 23385 6403 23443 6409
rect 23937 6443 23995 6449
rect 23937 6409 23949 6443
rect 23983 6440 23995 6443
rect 23983 6412 27476 6440
rect 23983 6409 23995 6412
rect 23937 6403 23995 6409
rect 9631 6344 12664 6372
rect 9631 6341 9643 6344
rect 9585 6335 9643 6341
rect 13354 6332 13360 6384
rect 13412 6372 13418 6384
rect 13412 6344 13768 6372
rect 13412 6332 13418 6344
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 992 6276 1593 6304
rect 992 6264 998 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 1581 6267 1639 6273
rect 2700 6276 2789 6304
rect 2700 6248 2728 6276
rect 2777 6273 2789 6276
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 2682 6196 2688 6248
rect 2740 6196 2746 6248
rect 2866 6196 2872 6248
rect 2924 6196 2930 6248
rect 3694 6236 3700 6248
rect 2976 6208 3700 6236
rect 1578 6128 1584 6180
rect 1636 6168 1642 6180
rect 2976 6168 3004 6208
rect 3694 6196 3700 6208
rect 3752 6196 3758 6248
rect 4062 6236 4068 6248
rect 3804 6208 4068 6236
rect 1636 6140 3004 6168
rect 1636 6128 1642 6140
rect 3418 6128 3424 6180
rect 3476 6168 3482 6180
rect 3804 6168 3832 6208
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 6380 6236 6408 6264
rect 6564 6236 6592 6267
rect 6380 6208 6592 6236
rect 6840 6236 6868 6267
rect 6914 6264 6920 6316
rect 6972 6264 6978 6316
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7550 6307 7608 6313
rect 7550 6304 7562 6307
rect 7156 6276 7562 6304
rect 7156 6264 7162 6276
rect 7550 6273 7562 6276
rect 7596 6273 7608 6307
rect 7550 6267 7608 6273
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 9180 6276 10793 6304
rect 9180 6264 9186 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 10962 6264 10968 6316
rect 11020 6264 11026 6316
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 11238 6304 11244 6316
rect 11195 6276 11244 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11238 6264 11244 6276
rect 11296 6304 11302 6316
rect 12710 6304 12716 6316
rect 11296 6276 12716 6304
rect 11296 6264 11302 6276
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 13740 6304 13768 6344
rect 13814 6332 13820 6384
rect 13872 6372 13878 6384
rect 15102 6372 15108 6384
rect 13872 6344 15108 6372
rect 13872 6332 13878 6344
rect 14568 6313 14596 6344
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 15838 6332 15844 6384
rect 15896 6332 15902 6384
rect 18506 6332 18512 6384
rect 18564 6332 18570 6384
rect 19794 6372 19800 6384
rect 19734 6344 19800 6372
rect 19794 6332 19800 6344
rect 19852 6332 19858 6384
rect 20254 6332 20260 6384
rect 20312 6372 20318 6384
rect 20622 6372 20628 6384
rect 20312 6344 20628 6372
rect 20312 6332 20318 6344
rect 20622 6332 20628 6344
rect 20680 6332 20686 6384
rect 20806 6332 20812 6384
rect 20864 6332 20870 6384
rect 23290 6372 23296 6384
rect 20916 6344 23296 6372
rect 14553 6307 14611 6313
rect 13740 6276 13952 6304
rect 13924 6248 13952 6276
rect 14553 6273 14565 6307
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6304 17187 6307
rect 17494 6304 17500 6316
rect 17175 6276 17500 6304
rect 17175 6273 17187 6276
rect 17129 6267 17187 6273
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 20916 6304 20944 6344
rect 23290 6332 23296 6344
rect 23348 6332 23354 6384
rect 24210 6332 24216 6384
rect 24268 6372 24274 6384
rect 24305 6375 24363 6381
rect 24305 6372 24317 6375
rect 24268 6344 24317 6372
rect 24268 6332 24274 6344
rect 24305 6341 24317 6344
rect 24351 6341 24363 6375
rect 24305 6335 24363 6341
rect 24397 6375 24455 6381
rect 24397 6341 24409 6375
rect 24443 6372 24455 6375
rect 24762 6372 24768 6384
rect 24443 6344 24768 6372
rect 24443 6341 24455 6344
rect 24397 6335 24455 6341
rect 24762 6332 24768 6344
rect 24820 6332 24826 6384
rect 25498 6332 25504 6384
rect 25556 6332 25562 6384
rect 27448 6381 27476 6412
rect 27522 6400 27528 6452
rect 27580 6440 27586 6452
rect 30282 6440 30288 6452
rect 27580 6412 30288 6440
rect 27580 6400 27586 6412
rect 30282 6400 30288 6412
rect 30340 6400 30346 6452
rect 31754 6400 31760 6452
rect 31812 6440 31818 6452
rect 31812 6412 32812 6440
rect 31812 6400 31818 6412
rect 27433 6375 27491 6381
rect 27433 6341 27445 6375
rect 27479 6341 27491 6375
rect 27433 6335 27491 6341
rect 27890 6332 27896 6384
rect 27948 6332 27954 6384
rect 29914 6372 29920 6384
rect 28736 6344 29920 6372
rect 19720 6276 20944 6304
rect 19720 6248 19748 6276
rect 22094 6264 22100 6316
rect 22152 6304 22158 6316
rect 22152 6276 22692 6304
rect 22152 6264 22158 6276
rect 7006 6236 7012 6248
rect 6840 6208 7012 6236
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 12805 6239 12863 6245
rect 7883 6208 12204 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 7558 6168 7564 6180
rect 3476 6140 3832 6168
rect 5368 6140 7564 6168
rect 3476 6128 3482 6140
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 2317 6103 2375 6109
rect 2317 6100 2329 6103
rect 1912 6072 2329 6100
rect 1912 6060 1918 6072
rect 2317 6069 2329 6072
rect 2363 6069 2375 6103
rect 2317 6063 2375 6069
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 5368 6100 5396 6140
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 12066 6168 12072 6180
rect 9364 6140 12072 6168
rect 9364 6128 9370 6140
rect 12066 6128 12072 6140
rect 12124 6128 12130 6180
rect 12176 6177 12204 6208
rect 12805 6205 12817 6239
rect 12851 6236 12863 6239
rect 13078 6236 13084 6248
rect 12851 6208 13084 6236
rect 12851 6205 12863 6208
rect 12805 6199 12863 6205
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 12161 6171 12219 6177
rect 12161 6137 12173 6171
rect 12207 6137 12219 6171
rect 13832 6168 13860 6199
rect 13906 6196 13912 6248
rect 13964 6196 13970 6248
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 14829 6239 14887 6245
rect 14829 6236 14841 6239
rect 14516 6208 14841 6236
rect 14516 6196 14522 6208
rect 14829 6205 14841 6208
rect 14875 6205 14887 6239
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 14829 6199 14887 6205
rect 15856 6208 17417 6236
rect 14550 6168 14556 6180
rect 13832 6140 14556 6168
rect 12161 6131 12219 6137
rect 14550 6128 14556 6140
rect 14608 6128 14614 6180
rect 4580 6072 5396 6100
rect 4580 6060 4586 6072
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 10413 6103 10471 6109
rect 10413 6100 10425 6103
rect 5500 6072 10425 6100
rect 5500 6060 5506 6072
rect 10413 6069 10425 6072
rect 10459 6069 10471 6103
rect 10413 6063 10471 6069
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 10689 6103 10747 6109
rect 10689 6100 10701 6103
rect 10560 6072 10701 6100
rect 10560 6060 10566 6072
rect 10689 6069 10701 6072
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 10778 6060 10784 6112
rect 10836 6100 10842 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10836 6072 10885 6100
rect 10836 6060 10842 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 10873 6063 10931 6069
rect 13354 6060 13360 6112
rect 13412 6060 13418 6112
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 15856 6100 15884 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18233 6239 18291 6245
rect 18233 6236 18245 6239
rect 17920 6208 18245 6236
rect 17920 6196 17926 6208
rect 18233 6205 18245 6208
rect 18279 6205 18291 6239
rect 18966 6236 18972 6248
rect 18233 6199 18291 6205
rect 18340 6208 18972 6236
rect 16022 6128 16028 6180
rect 16080 6168 16086 6180
rect 16301 6171 16359 6177
rect 16301 6168 16313 6171
rect 16080 6140 16313 6168
rect 16080 6128 16086 6140
rect 16301 6137 16313 6140
rect 16347 6168 16359 6171
rect 18340 6168 18368 6208
rect 18966 6196 18972 6208
rect 19024 6196 19030 6248
rect 19702 6196 19708 6248
rect 19760 6196 19766 6248
rect 19981 6239 20039 6245
rect 19981 6205 19993 6239
rect 20027 6236 20039 6239
rect 20346 6236 20352 6248
rect 20027 6208 20352 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 20346 6196 20352 6208
rect 20404 6196 20410 6248
rect 20806 6196 20812 6248
rect 20864 6236 20870 6248
rect 20901 6239 20959 6245
rect 20901 6236 20913 6239
rect 20864 6208 20913 6236
rect 20864 6196 20870 6208
rect 20901 6205 20913 6208
rect 20947 6205 20959 6239
rect 20901 6199 20959 6205
rect 21085 6239 21143 6245
rect 21085 6205 21097 6239
rect 21131 6236 21143 6239
rect 22278 6236 22284 6248
rect 21131 6208 22284 6236
rect 21131 6205 21143 6208
rect 21085 6199 21143 6205
rect 20441 6171 20499 6177
rect 20441 6168 20453 6171
rect 16347 6140 18368 6168
rect 19536 6140 20453 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 13688 6072 15884 6100
rect 13688 6060 13694 6072
rect 16574 6060 16580 6112
rect 16632 6100 16638 6112
rect 19536 6100 19564 6140
rect 20441 6137 20453 6140
rect 20487 6137 20499 6171
rect 20441 6131 20499 6137
rect 20530 6128 20536 6180
rect 20588 6168 20594 6180
rect 21100 6168 21128 6199
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 22373 6239 22431 6245
rect 22373 6205 22385 6239
rect 22419 6205 22431 6239
rect 22664 6236 22692 6276
rect 22738 6264 22744 6316
rect 22796 6304 22802 6316
rect 23201 6307 23259 6313
rect 23201 6304 23213 6307
rect 22796 6276 23213 6304
rect 22796 6264 22802 6276
rect 23201 6273 23213 6276
rect 23247 6273 23259 6307
rect 25774 6304 25780 6316
rect 23201 6267 23259 6273
rect 23676 6276 25780 6304
rect 23566 6236 23572 6248
rect 22664 6208 23572 6236
rect 22373 6199 22431 6205
rect 20588 6140 21128 6168
rect 20588 6128 20594 6140
rect 22094 6128 22100 6180
rect 22152 6168 22158 6180
rect 22388 6168 22416 6199
rect 23566 6196 23572 6208
rect 23624 6196 23630 6248
rect 22152 6140 22416 6168
rect 22152 6128 22158 6140
rect 23014 6128 23020 6180
rect 23072 6168 23078 6180
rect 23676 6168 23704 6276
rect 24596 6245 24624 6276
rect 25774 6264 25780 6276
rect 25832 6304 25838 6316
rect 26142 6304 26148 6316
rect 25832 6276 26148 6304
rect 25832 6264 25838 6276
rect 26142 6264 26148 6276
rect 26200 6264 26206 6316
rect 24581 6239 24639 6245
rect 24581 6205 24593 6239
rect 24627 6205 24639 6239
rect 24581 6199 24639 6205
rect 25130 6196 25136 6248
rect 25188 6236 25194 6248
rect 26329 6239 26387 6245
rect 26329 6236 26341 6239
rect 25188 6208 26341 6236
rect 25188 6196 25194 6208
rect 26329 6205 26341 6208
rect 26375 6236 26387 6239
rect 27157 6239 27215 6245
rect 27157 6236 27169 6239
rect 26375 6208 27169 6236
rect 26375 6205 26387 6208
rect 26329 6199 26387 6205
rect 27157 6205 27169 6208
rect 27203 6205 27215 6239
rect 28736 6236 28764 6344
rect 29914 6332 29920 6344
rect 29972 6332 29978 6384
rect 31386 6372 31392 6384
rect 31142 6344 31392 6372
rect 31386 6332 31392 6344
rect 31444 6332 31450 6384
rect 32674 6332 32680 6384
rect 32732 6332 32738 6384
rect 32784 6372 32812 6412
rect 33704 6412 34008 6440
rect 33704 6372 33732 6412
rect 32784 6344 33732 6372
rect 33781 6375 33839 6381
rect 31294 6264 31300 6316
rect 31352 6304 31358 6316
rect 32490 6304 32496 6316
rect 31352 6276 32496 6304
rect 31352 6264 31358 6276
rect 32490 6264 32496 6276
rect 32548 6304 32554 6316
rect 33658 6313 33686 6344
rect 33781 6341 33793 6375
rect 33827 6341 33839 6375
rect 33781 6335 33839 6341
rect 33643 6307 33701 6313
rect 32548 6276 33548 6304
rect 32548 6264 32554 6276
rect 27157 6199 27215 6205
rect 27264 6208 28764 6236
rect 23072 6140 23704 6168
rect 23072 6128 23078 6140
rect 26510 6128 26516 6180
rect 26568 6168 26574 6180
rect 27264 6168 27292 6208
rect 29362 6196 29368 6248
rect 29420 6236 29426 6248
rect 29641 6239 29699 6245
rect 29641 6236 29653 6239
rect 29420 6208 29653 6236
rect 29420 6196 29426 6208
rect 29641 6205 29653 6208
rect 29687 6205 29699 6239
rect 29641 6199 29699 6205
rect 29917 6239 29975 6245
rect 29917 6205 29929 6239
rect 29963 6236 29975 6239
rect 29963 6208 31754 6236
rect 29963 6205 29975 6208
rect 29917 6199 29975 6205
rect 26568 6140 27292 6168
rect 31726 6168 31754 6208
rect 32674 6196 32680 6248
rect 32732 6236 32738 6248
rect 32769 6239 32827 6245
rect 32769 6236 32781 6239
rect 32732 6208 32781 6236
rect 32732 6196 32738 6208
rect 32769 6205 32781 6208
rect 32815 6205 32827 6239
rect 32769 6199 32827 6205
rect 32953 6239 33011 6245
rect 32953 6205 32965 6239
rect 32999 6236 33011 6239
rect 33042 6236 33048 6248
rect 32999 6208 33048 6236
rect 32999 6205 33011 6208
rect 32953 6199 33011 6205
rect 33042 6196 33048 6208
rect 33100 6196 33106 6248
rect 33520 6236 33548 6276
rect 33643 6273 33655 6307
rect 33689 6273 33701 6307
rect 33643 6267 33701 6273
rect 33796 6236 33824 6335
rect 33870 6332 33876 6384
rect 33928 6332 33934 6384
rect 33980 6372 34008 6412
rect 34146 6400 34152 6452
rect 34204 6400 34210 6452
rect 36357 6443 36415 6449
rect 36357 6440 36369 6443
rect 34256 6412 36369 6440
rect 34256 6372 34284 6412
rect 36357 6409 36369 6412
rect 36403 6409 36415 6443
rect 36357 6403 36415 6409
rect 37090 6400 37096 6452
rect 37148 6440 37154 6452
rect 37461 6443 37519 6449
rect 37461 6440 37473 6443
rect 37148 6412 37473 6440
rect 37148 6400 37154 6412
rect 37461 6409 37473 6412
rect 37507 6409 37519 6443
rect 37461 6403 37519 6409
rect 37921 6443 37979 6449
rect 37921 6409 37933 6443
rect 37967 6440 37979 6443
rect 38470 6440 38476 6452
rect 37967 6412 38476 6440
rect 37967 6409 37979 6412
rect 37921 6403 37979 6409
rect 38470 6400 38476 6412
rect 38528 6400 38534 6452
rect 36538 6372 36544 6384
rect 33980 6344 34284 6372
rect 36110 6344 36544 6372
rect 36538 6332 36544 6344
rect 36596 6332 36602 6384
rect 33962 6264 33968 6316
rect 34020 6264 34026 6316
rect 36170 6264 36176 6316
rect 36228 6304 36234 6316
rect 37829 6307 37887 6313
rect 37829 6304 37841 6307
rect 36228 6276 37841 6304
rect 36228 6264 36234 6276
rect 37829 6273 37841 6276
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 33520 6208 33824 6236
rect 34238 6196 34244 6248
rect 34296 6236 34302 6248
rect 34609 6239 34667 6245
rect 34609 6236 34621 6239
rect 34296 6208 34621 6236
rect 34296 6196 34302 6208
rect 34609 6205 34621 6208
rect 34655 6236 34667 6239
rect 34655 6208 34744 6236
rect 34655 6205 34667 6208
rect 34609 6199 34667 6205
rect 32309 6171 32367 6177
rect 32309 6168 32321 6171
rect 31726 6140 32321 6168
rect 26568 6128 26574 6140
rect 32309 6137 32321 6140
rect 32355 6137 32367 6171
rect 32309 6131 32367 6137
rect 16632 6072 19564 6100
rect 16632 6060 16638 6072
rect 19886 6060 19892 6112
rect 19944 6100 19950 6112
rect 22186 6100 22192 6112
rect 19944 6072 22192 6100
rect 19944 6060 19950 6072
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 24762 6060 24768 6112
rect 24820 6100 24826 6112
rect 26234 6100 26240 6112
rect 24820 6072 26240 6100
rect 24820 6060 24826 6072
rect 26234 6060 26240 6072
rect 26292 6100 26298 6112
rect 28905 6103 28963 6109
rect 28905 6100 28917 6103
rect 26292 6072 28917 6100
rect 26292 6060 26298 6072
rect 28905 6069 28917 6072
rect 28951 6069 28963 6103
rect 28905 6063 28963 6069
rect 29086 6060 29092 6112
rect 29144 6100 29150 6112
rect 30098 6100 30104 6112
rect 29144 6072 30104 6100
rect 29144 6060 29150 6072
rect 30098 6060 30104 6072
rect 30156 6060 30162 6112
rect 31294 6060 31300 6112
rect 31352 6100 31358 6112
rect 31389 6103 31447 6109
rect 31389 6100 31401 6103
rect 31352 6072 31401 6100
rect 31352 6060 31358 6072
rect 31389 6069 31401 6072
rect 31435 6100 31447 6103
rect 32674 6100 32680 6112
rect 31435 6072 32680 6100
rect 31435 6069 31447 6072
rect 31389 6063 31447 6069
rect 32674 6060 32680 6072
rect 32732 6060 32738 6112
rect 32766 6060 32772 6112
rect 32824 6100 32830 6112
rect 34146 6100 34152 6112
rect 32824 6072 34152 6100
rect 32824 6060 32830 6072
rect 34146 6060 34152 6072
rect 34204 6060 34210 6112
rect 34716 6100 34744 6208
rect 34882 6196 34888 6248
rect 34940 6196 34946 6248
rect 35618 6196 35624 6248
rect 35676 6236 35682 6248
rect 37918 6236 37924 6248
rect 35676 6208 37924 6236
rect 35676 6196 35682 6208
rect 37918 6196 37924 6208
rect 37976 6196 37982 6248
rect 38013 6239 38071 6245
rect 38013 6205 38025 6239
rect 38059 6205 38071 6239
rect 38013 6199 38071 6205
rect 35986 6128 35992 6180
rect 36044 6168 36050 6180
rect 38028 6168 38056 6199
rect 36044 6140 38056 6168
rect 36044 6128 36050 6140
rect 35894 6100 35900 6112
rect 34716 6072 35900 6100
rect 35894 6060 35900 6072
rect 35952 6060 35958 6112
rect 1104 6010 39192 6032
rect 1104 5958 5711 6010
rect 5763 5958 5775 6010
rect 5827 5958 5839 6010
rect 5891 5958 5903 6010
rect 5955 5958 5967 6010
rect 6019 5958 15233 6010
rect 15285 5958 15297 6010
rect 15349 5958 15361 6010
rect 15413 5958 15425 6010
rect 15477 5958 15489 6010
rect 15541 5958 24755 6010
rect 24807 5958 24819 6010
rect 24871 5958 24883 6010
rect 24935 5958 24947 6010
rect 24999 5958 25011 6010
rect 25063 5958 34277 6010
rect 34329 5958 34341 6010
rect 34393 5958 34405 6010
rect 34457 5958 34469 6010
rect 34521 5958 34533 6010
rect 34585 5958 39192 6010
rect 1104 5936 39192 5958
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 2004 5868 3648 5896
rect 2004 5856 2010 5868
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2314 5760 2320 5772
rect 1995 5732 2320 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 2314 5720 2320 5732
rect 2372 5720 2378 5772
rect 1578 5652 1584 5704
rect 1636 5692 1642 5704
rect 1673 5695 1731 5701
rect 1673 5692 1685 5695
rect 1636 5664 1685 5692
rect 1636 5652 1642 5664
rect 1673 5661 1685 5664
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 3234 5624 3240 5636
rect 3174 5596 3240 5624
rect 3234 5584 3240 5596
rect 3292 5584 3298 5636
rect 3620 5624 3648 5868
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 7082 5899 7140 5905
rect 7082 5896 7094 5899
rect 5316 5868 7094 5896
rect 5316 5856 5322 5868
rect 7082 5865 7094 5868
rect 7128 5865 7140 5899
rect 7082 5859 7140 5865
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 8294 5896 8300 5908
rect 7616 5868 8300 5896
rect 7616 5856 7622 5868
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 8846 5896 8852 5908
rect 8619 5868 8852 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 8956 5868 10456 5896
rect 6270 5788 6276 5840
rect 6328 5828 6334 5840
rect 6822 5828 6828 5840
rect 6328 5800 6828 5828
rect 6328 5788 6334 5800
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8956 5828 8984 5868
rect 8168 5800 8984 5828
rect 10428 5828 10456 5868
rect 10870 5856 10876 5908
rect 10928 5856 10934 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 13722 5896 13728 5908
rect 13044 5868 13728 5896
rect 13044 5856 13050 5868
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 14458 5856 14464 5908
rect 14516 5856 14522 5908
rect 14550 5856 14556 5908
rect 14608 5896 14614 5908
rect 15746 5896 15752 5908
rect 14608 5868 15752 5896
rect 14608 5856 14614 5868
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 17770 5856 17776 5908
rect 17828 5896 17834 5908
rect 19429 5899 19487 5905
rect 19429 5896 19441 5899
rect 17828 5868 19441 5896
rect 17828 5856 17834 5868
rect 19429 5865 19441 5868
rect 19475 5865 19487 5899
rect 19429 5859 19487 5865
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 20622 5896 20628 5908
rect 19668 5868 20628 5896
rect 19668 5856 19674 5868
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 23014 5896 23020 5908
rect 20916 5868 23020 5896
rect 11974 5828 11980 5840
rect 10428 5800 11980 5828
rect 8168 5788 8174 5800
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 14826 5788 14832 5840
rect 14884 5828 14890 5840
rect 14884 5800 15056 5828
rect 14884 5788 14890 5800
rect 3694 5720 3700 5772
rect 3752 5760 3758 5772
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 3752 5732 4629 5760
rect 3752 5720 3758 5732
rect 4617 5729 4629 5732
rect 4663 5760 4675 5763
rect 8386 5760 8392 5772
rect 4663 5732 6592 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 6564 5704 6592 5732
rect 6840 5732 8392 5760
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4522 5692 4528 5704
rect 4019 5664 4528 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 6546 5652 6552 5704
rect 6604 5692 6610 5704
rect 6840 5701 6868 5732
rect 8386 5720 8392 5732
rect 8444 5760 8450 5772
rect 9125 5763 9183 5769
rect 9125 5760 9137 5763
rect 8444 5732 9137 5760
rect 8444 5720 8450 5732
rect 9125 5729 9137 5732
rect 9171 5729 9183 5763
rect 9125 5723 9183 5729
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5760 9459 5763
rect 11054 5760 11060 5772
rect 9447 5732 11060 5760
rect 9447 5729 9459 5732
rect 9401 5723 9459 5729
rect 11054 5720 11060 5732
rect 11112 5720 11118 5772
rect 12253 5763 12311 5769
rect 12253 5729 12265 5763
rect 12299 5760 12311 5763
rect 12299 5732 13768 5760
rect 12299 5729 12311 5732
rect 12253 5723 12311 5729
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6604 5664 6837 5692
rect 6604 5652 6610 5664
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 11388 5664 11989 5692
rect 11388 5652 11394 5664
rect 11977 5661 11989 5664
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 3620 5596 4844 5624
rect 3421 5559 3479 5565
rect 3421 5525 3433 5559
rect 3467 5556 3479 5559
rect 3970 5556 3976 5568
rect 3467 5528 3976 5556
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4062 5516 4068 5568
rect 4120 5516 4126 5568
rect 4816 5556 4844 5596
rect 4890 5584 4896 5636
rect 4948 5584 4954 5636
rect 6178 5624 6184 5636
rect 6118 5596 6184 5624
rect 6178 5584 6184 5596
rect 6236 5584 6242 5636
rect 6638 5584 6644 5636
rect 6696 5624 6702 5636
rect 11790 5624 11796 5636
rect 6696 5596 7590 5624
rect 10626 5596 11796 5624
rect 6696 5584 6702 5596
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 13538 5624 13544 5636
rect 13478 5596 13544 5624
rect 13538 5584 13544 5596
rect 13596 5584 13602 5636
rect 13740 5624 13768 5732
rect 14918 5720 14924 5772
rect 14976 5720 14982 5772
rect 15028 5769 15056 5800
rect 18138 5788 18144 5840
rect 18196 5788 18202 5840
rect 19702 5828 19708 5840
rect 18616 5800 19708 5828
rect 15013 5763 15071 5769
rect 15013 5729 15025 5763
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 15930 5720 15936 5772
rect 15988 5720 15994 5772
rect 17405 5763 17463 5769
rect 17405 5729 17417 5763
rect 17451 5760 17463 5763
rect 18616 5760 18644 5800
rect 19702 5788 19708 5800
rect 19760 5788 19766 5840
rect 19797 5831 19855 5837
rect 19797 5797 19809 5831
rect 19843 5828 19855 5831
rect 20806 5828 20812 5840
rect 19843 5800 20812 5828
rect 19843 5797 19855 5800
rect 19797 5791 19855 5797
rect 20806 5788 20812 5800
rect 20864 5788 20870 5840
rect 17451 5732 18644 5760
rect 17451 5729 17463 5732
rect 17405 5723 17463 5729
rect 18690 5720 18696 5772
rect 18748 5760 18754 5772
rect 19886 5760 19892 5772
rect 18748 5732 19892 5760
rect 18748 5720 18754 5732
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 20916 5769 20944 5868
rect 23014 5856 23020 5868
rect 23072 5856 23078 5908
rect 23198 5856 23204 5908
rect 23256 5856 23262 5908
rect 23845 5899 23903 5905
rect 23845 5865 23857 5899
rect 23891 5896 23903 5899
rect 24578 5896 24584 5908
rect 23891 5868 24584 5896
rect 23891 5865 23903 5868
rect 23845 5859 23903 5865
rect 24578 5856 24584 5868
rect 24636 5856 24642 5908
rect 25133 5899 25191 5905
rect 25133 5865 25145 5899
rect 25179 5896 25191 5899
rect 25406 5896 25412 5908
rect 25179 5868 25412 5896
rect 25179 5865 25191 5868
rect 25133 5859 25191 5865
rect 25406 5856 25412 5868
rect 25464 5856 25470 5908
rect 26326 5856 26332 5908
rect 26384 5896 26390 5908
rect 26881 5899 26939 5905
rect 26881 5896 26893 5899
rect 26384 5868 26893 5896
rect 26384 5856 26390 5868
rect 26881 5865 26893 5868
rect 26927 5865 26939 5899
rect 30929 5899 30987 5905
rect 26881 5859 26939 5865
rect 27080 5868 30880 5896
rect 24029 5831 24087 5837
rect 24029 5797 24041 5831
rect 24075 5828 24087 5831
rect 26050 5828 26056 5840
rect 24075 5800 26056 5828
rect 24075 5797 24087 5800
rect 24029 5791 24087 5797
rect 26050 5788 26056 5800
rect 26108 5788 26114 5840
rect 26418 5788 26424 5840
rect 26476 5828 26482 5840
rect 26513 5831 26571 5837
rect 26513 5828 26525 5831
rect 26476 5800 26525 5828
rect 26476 5788 26482 5800
rect 26513 5797 26525 5800
rect 26559 5797 26571 5831
rect 26513 5791 26571 5797
rect 27080 5772 27108 5868
rect 27709 5831 27767 5837
rect 27709 5797 27721 5831
rect 27755 5828 27767 5831
rect 30006 5828 30012 5840
rect 27755 5800 30012 5828
rect 27755 5797 27767 5800
rect 27709 5791 27767 5797
rect 30006 5788 30012 5800
rect 30064 5788 30070 5840
rect 30098 5788 30104 5840
rect 30156 5828 30162 5840
rect 30742 5828 30748 5840
rect 30156 5800 30748 5828
rect 30156 5788 30162 5800
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 21453 5763 21511 5769
rect 21453 5729 21465 5763
rect 21499 5760 21511 5763
rect 25130 5760 25136 5772
rect 21499 5732 25136 5760
rect 21499 5729 21511 5732
rect 21453 5723 21511 5729
rect 25130 5720 25136 5732
rect 25188 5720 25194 5772
rect 25590 5760 25596 5772
rect 25240 5732 25596 5760
rect 14090 5652 14096 5704
rect 14148 5692 14154 5704
rect 14550 5692 14556 5704
rect 14148 5664 14556 5692
rect 14148 5652 14154 5664
rect 14550 5652 14556 5664
rect 14608 5652 14614 5704
rect 15470 5692 15476 5704
rect 14844 5664 15476 5692
rect 14844 5624 14872 5664
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 15654 5652 15660 5704
rect 15712 5652 15718 5704
rect 17310 5692 17316 5704
rect 17066 5664 17316 5692
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 18322 5652 18328 5704
rect 18380 5692 18386 5704
rect 18601 5695 18659 5701
rect 18601 5692 18613 5695
rect 18380 5664 18613 5692
rect 18380 5652 18386 5664
rect 18601 5661 18613 5664
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 19392 5664 19441 5692
rect 19392 5652 19398 5664
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 19429 5655 19487 5661
rect 19610 5652 19616 5704
rect 19668 5652 19674 5704
rect 20622 5652 20628 5704
rect 20680 5652 20686 5704
rect 20717 5695 20775 5701
rect 20717 5661 20729 5695
rect 20763 5692 20775 5695
rect 21082 5692 21088 5704
rect 20763 5664 21088 5692
rect 20763 5661 20775 5664
rect 20717 5655 20775 5661
rect 21082 5652 21088 5664
rect 21140 5652 21146 5704
rect 24857 5695 24915 5701
rect 24857 5692 24869 5695
rect 23032 5664 24869 5692
rect 16022 5624 16028 5636
rect 13740 5596 14872 5624
rect 15396 5596 16028 5624
rect 5166 5556 5172 5568
rect 4816 5528 5172 5556
rect 5166 5516 5172 5528
rect 5224 5556 5230 5568
rect 6365 5559 6423 5565
rect 6365 5556 6377 5559
rect 5224 5528 6377 5556
rect 5224 5516 5230 5528
rect 6365 5525 6377 5528
rect 6411 5525 6423 5559
rect 6365 5519 6423 5525
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 11422 5556 11428 5568
rect 9824 5528 11428 5556
rect 9824 5516 9830 5528
rect 11422 5516 11428 5528
rect 11480 5556 11486 5568
rect 12066 5556 12072 5568
rect 11480 5528 12072 5556
rect 11480 5516 11486 5528
rect 12066 5516 12072 5528
rect 12124 5556 12130 5568
rect 13630 5556 13636 5568
rect 12124 5528 13636 5556
rect 12124 5516 12130 5528
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 13725 5559 13783 5565
rect 13725 5525 13737 5559
rect 13771 5556 13783 5559
rect 14734 5556 14740 5568
rect 13771 5528 14740 5556
rect 13771 5525 13783 5528
rect 13725 5519 13783 5525
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 14829 5559 14887 5565
rect 14829 5525 14841 5559
rect 14875 5556 14887 5559
rect 15396 5556 15424 5596
rect 16022 5584 16028 5596
rect 16080 5584 16086 5636
rect 20640 5624 20668 5652
rect 21174 5624 21180 5636
rect 17236 5596 20300 5624
rect 20640 5596 21180 5624
rect 14875 5528 15424 5556
rect 14875 5525 14887 5528
rect 14829 5519 14887 5525
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 17236 5556 17264 5596
rect 15528 5528 17264 5556
rect 15528 5516 15534 5528
rect 17310 5516 17316 5568
rect 17368 5556 17374 5568
rect 17954 5556 17960 5568
rect 17368 5528 17960 5556
rect 17368 5516 17374 5528
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 18509 5559 18567 5565
rect 18509 5525 18521 5559
rect 18555 5556 18567 5559
rect 19058 5556 19064 5568
rect 18555 5528 19064 5556
rect 18555 5525 18567 5528
rect 18509 5519 18567 5525
rect 19058 5516 19064 5528
rect 19116 5516 19122 5568
rect 20272 5565 20300 5596
rect 21174 5584 21180 5596
rect 21232 5584 21238 5636
rect 21634 5584 21640 5636
rect 21692 5624 21698 5636
rect 21729 5627 21787 5633
rect 21729 5624 21741 5627
rect 21692 5596 21741 5624
rect 21692 5584 21698 5596
rect 21729 5593 21741 5596
rect 21775 5593 21787 5627
rect 21729 5587 21787 5593
rect 22370 5584 22376 5636
rect 22428 5584 22434 5636
rect 20257 5559 20315 5565
rect 20257 5525 20269 5559
rect 20303 5525 20315 5559
rect 20257 5519 20315 5525
rect 22554 5516 22560 5568
rect 22612 5556 22618 5568
rect 23032 5556 23060 5664
rect 24857 5661 24869 5664
rect 24903 5692 24915 5695
rect 25240 5692 25268 5732
rect 25590 5720 25596 5732
rect 25648 5720 25654 5772
rect 25777 5763 25835 5769
rect 25777 5729 25789 5763
rect 25823 5760 25835 5763
rect 25958 5760 25964 5772
rect 25823 5732 25964 5760
rect 25823 5729 25835 5732
rect 25777 5723 25835 5729
rect 25958 5720 25964 5732
rect 26016 5720 26022 5772
rect 26878 5720 26884 5772
rect 26936 5760 26942 5772
rect 26973 5763 27031 5769
rect 26973 5760 26985 5763
rect 26936 5732 26985 5760
rect 26936 5720 26942 5732
rect 26973 5729 26985 5732
rect 27019 5729 27031 5763
rect 26973 5723 27031 5729
rect 27062 5720 27068 5772
rect 27120 5720 27126 5772
rect 27798 5720 27804 5772
rect 27856 5760 27862 5772
rect 28169 5763 28227 5769
rect 28169 5760 28181 5763
rect 27856 5732 28181 5760
rect 27856 5720 27862 5732
rect 28169 5729 28181 5732
rect 28215 5729 28227 5763
rect 28169 5723 28227 5729
rect 28353 5763 28411 5769
rect 28353 5729 28365 5763
rect 28399 5729 28411 5763
rect 28353 5723 28411 5729
rect 24903 5664 25268 5692
rect 24903 5661 24915 5664
rect 24857 5655 24915 5661
rect 25314 5652 25320 5704
rect 25372 5692 25378 5704
rect 25501 5695 25559 5701
rect 25501 5692 25513 5695
rect 25372 5664 25513 5692
rect 25372 5652 25378 5664
rect 25501 5661 25513 5664
rect 25547 5661 25559 5695
rect 25501 5655 25559 5661
rect 26786 5652 26792 5704
rect 26844 5652 26850 5704
rect 27249 5695 27307 5701
rect 27249 5661 27261 5695
rect 27295 5692 27307 5695
rect 27430 5692 27436 5704
rect 27295 5664 27436 5692
rect 27295 5661 27307 5664
rect 27249 5655 27307 5661
rect 27430 5652 27436 5664
rect 27488 5652 27494 5704
rect 27614 5652 27620 5704
rect 27672 5692 27678 5704
rect 27982 5692 27988 5704
rect 27672 5664 27988 5692
rect 27672 5652 27678 5664
rect 27982 5652 27988 5664
rect 28040 5652 28046 5704
rect 28074 5652 28080 5704
rect 28132 5652 28138 5704
rect 23661 5627 23719 5633
rect 23661 5593 23673 5627
rect 23707 5624 23719 5627
rect 24762 5624 24768 5636
rect 23707 5596 24768 5624
rect 23707 5593 23719 5596
rect 23661 5587 23719 5593
rect 24762 5584 24768 5596
rect 24820 5584 24826 5636
rect 26694 5584 26700 5636
rect 26752 5624 26758 5636
rect 27522 5624 27528 5636
rect 26752 5596 27528 5624
rect 26752 5584 26758 5596
rect 27522 5584 27528 5596
rect 27580 5584 27586 5636
rect 28368 5624 28396 5723
rect 28534 5720 28540 5772
rect 28592 5760 28598 5772
rect 29914 5760 29920 5772
rect 28592 5732 29920 5760
rect 28592 5720 28598 5732
rect 29914 5720 29920 5732
rect 29972 5720 29978 5772
rect 30300 5769 30328 5800
rect 30742 5788 30748 5800
rect 30800 5788 30806 5840
rect 30852 5828 30880 5868
rect 30929 5865 30941 5899
rect 30975 5896 30987 5899
rect 34882 5896 34888 5908
rect 30975 5868 34888 5896
rect 30975 5865 30987 5868
rect 30929 5859 30987 5865
rect 34882 5856 34888 5868
rect 34940 5856 34946 5908
rect 35342 5856 35348 5908
rect 35400 5896 35406 5908
rect 35400 5868 37964 5896
rect 35400 5856 35406 5868
rect 32398 5828 32404 5840
rect 30852 5800 32404 5828
rect 32398 5788 32404 5800
rect 32456 5788 32462 5840
rect 30285 5763 30343 5769
rect 30285 5729 30297 5763
rect 30331 5729 30343 5763
rect 30285 5723 30343 5729
rect 30374 5720 30380 5772
rect 30432 5760 30438 5772
rect 30926 5760 30932 5772
rect 30432 5732 30932 5760
rect 30432 5720 30438 5732
rect 30926 5720 30932 5732
rect 30984 5760 30990 5772
rect 31481 5763 31539 5769
rect 31481 5760 31493 5763
rect 30984 5732 31493 5760
rect 30984 5720 30990 5732
rect 31481 5729 31493 5732
rect 31527 5729 31539 5763
rect 31481 5723 31539 5729
rect 32030 5720 32036 5772
rect 32088 5760 32094 5772
rect 32585 5763 32643 5769
rect 32585 5760 32597 5763
rect 32088 5732 32597 5760
rect 32088 5720 32094 5732
rect 32585 5729 32597 5732
rect 32631 5760 32643 5763
rect 33502 5760 33508 5772
rect 32631 5732 33508 5760
rect 32631 5729 32643 5732
rect 32585 5723 32643 5729
rect 33502 5720 33508 5732
rect 33560 5720 33566 5772
rect 33980 5732 35848 5760
rect 28442 5652 28448 5704
rect 28500 5692 28506 5704
rect 31294 5692 31300 5704
rect 28500 5664 31300 5692
rect 28500 5652 28506 5664
rect 31294 5652 31300 5664
rect 31352 5652 31358 5704
rect 31389 5695 31447 5701
rect 31389 5661 31401 5695
rect 31435 5692 31447 5695
rect 31754 5692 31760 5704
rect 31435 5664 31760 5692
rect 31435 5661 31447 5664
rect 31389 5655 31447 5661
rect 31754 5652 31760 5664
rect 31812 5652 31818 5704
rect 33980 5678 34008 5732
rect 34606 5652 34612 5704
rect 34664 5692 34670 5704
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 34664 5664 34897 5692
rect 34664 5652 34670 5664
rect 34885 5661 34897 5664
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 35069 5695 35127 5701
rect 35069 5661 35081 5695
rect 35115 5692 35127 5695
rect 35434 5692 35440 5704
rect 35115 5664 35440 5692
rect 35115 5661 35127 5664
rect 35069 5655 35127 5661
rect 35434 5652 35440 5664
rect 35492 5652 35498 5704
rect 28368 5596 28488 5624
rect 22612 5528 23060 5556
rect 23871 5559 23929 5565
rect 22612 5516 22618 5528
rect 23871 5525 23883 5559
rect 23917 5556 23929 5559
rect 25866 5556 25872 5568
rect 23917 5528 25872 5556
rect 23917 5525 23929 5528
rect 23871 5519 23929 5525
rect 25866 5516 25872 5528
rect 25924 5556 25930 5568
rect 27798 5556 27804 5568
rect 25924 5528 27804 5556
rect 25924 5516 25930 5528
rect 27798 5516 27804 5528
rect 27856 5516 27862 5568
rect 28460 5556 28488 5596
rect 28534 5584 28540 5636
rect 28592 5624 28598 5636
rect 28997 5627 29055 5633
rect 28997 5624 29009 5627
rect 28592 5596 29009 5624
rect 28592 5584 28598 5596
rect 28997 5593 29009 5596
rect 29043 5593 29055 5627
rect 28997 5587 29055 5593
rect 29270 5584 29276 5636
rect 29328 5624 29334 5636
rect 32861 5627 32919 5633
rect 29328 5596 31754 5624
rect 29328 5584 29334 5596
rect 28718 5556 28724 5568
rect 28460 5528 28724 5556
rect 28718 5516 28724 5528
rect 28776 5516 28782 5568
rect 29086 5516 29092 5568
rect 29144 5516 29150 5568
rect 29178 5516 29184 5568
rect 29236 5556 29242 5568
rect 29733 5559 29791 5565
rect 29733 5556 29745 5559
rect 29236 5528 29745 5556
rect 29236 5516 29242 5528
rect 29733 5525 29745 5528
rect 29779 5525 29791 5559
rect 29733 5519 29791 5525
rect 30098 5516 30104 5568
rect 30156 5516 30162 5568
rect 30193 5559 30251 5565
rect 30193 5525 30205 5559
rect 30239 5556 30251 5559
rect 30374 5556 30380 5568
rect 30239 5528 30380 5556
rect 30239 5525 30251 5528
rect 30193 5519 30251 5525
rect 30374 5516 30380 5528
rect 30432 5516 30438 5568
rect 30466 5516 30472 5568
rect 30524 5556 30530 5568
rect 31202 5556 31208 5568
rect 30524 5528 31208 5556
rect 30524 5516 30530 5528
rect 31202 5516 31208 5528
rect 31260 5556 31266 5568
rect 31297 5559 31355 5565
rect 31297 5556 31309 5559
rect 31260 5528 31309 5556
rect 31260 5516 31266 5528
rect 31297 5525 31309 5528
rect 31343 5525 31355 5559
rect 31726 5556 31754 5596
rect 32861 5593 32873 5627
rect 32907 5624 32919 5627
rect 32950 5624 32956 5636
rect 32907 5596 32956 5624
rect 32907 5593 32919 5596
rect 32861 5587 32919 5593
rect 32950 5584 32956 5596
rect 33008 5584 33014 5636
rect 35253 5627 35311 5633
rect 35253 5624 35265 5627
rect 34164 5596 35265 5624
rect 34164 5556 34192 5596
rect 35253 5593 35265 5596
rect 35299 5593 35311 5627
rect 35253 5587 35311 5593
rect 31726 5528 34192 5556
rect 31297 5519 31355 5525
rect 34238 5516 34244 5568
rect 34296 5556 34302 5568
rect 34333 5559 34391 5565
rect 34333 5556 34345 5559
rect 34296 5528 34345 5556
rect 34296 5516 34302 5528
rect 34333 5525 34345 5528
rect 34379 5556 34391 5559
rect 35618 5556 35624 5568
rect 34379 5528 35624 5556
rect 34379 5525 34391 5528
rect 34333 5519 34391 5525
rect 35618 5516 35624 5528
rect 35676 5516 35682 5568
rect 35820 5556 35848 5732
rect 35894 5720 35900 5772
rect 35952 5760 35958 5772
rect 36814 5760 36820 5772
rect 35952 5732 36820 5760
rect 35952 5720 35958 5732
rect 36814 5720 36820 5732
rect 36872 5720 36878 5772
rect 37936 5769 37964 5868
rect 38010 5856 38016 5908
rect 38068 5896 38074 5908
rect 38473 5899 38531 5905
rect 38473 5896 38485 5899
rect 38068 5868 38485 5896
rect 38068 5856 38074 5868
rect 38473 5865 38485 5868
rect 38519 5865 38531 5899
rect 38473 5859 38531 5865
rect 37921 5763 37979 5769
rect 37921 5729 37933 5763
rect 37967 5729 37979 5763
rect 37921 5723 37979 5729
rect 37274 5652 37280 5704
rect 37332 5652 37338 5704
rect 38378 5652 38384 5704
rect 38436 5652 38442 5704
rect 36078 5584 36084 5636
rect 36136 5624 36142 5636
rect 36173 5627 36231 5633
rect 36173 5624 36185 5627
rect 36136 5596 36185 5624
rect 36136 5584 36142 5596
rect 36173 5593 36185 5596
rect 36219 5593 36231 5627
rect 36173 5587 36231 5593
rect 37182 5556 37188 5568
rect 35820 5528 37188 5556
rect 37182 5516 37188 5528
rect 37240 5516 37246 5568
rect 1104 5466 39352 5488
rect 1104 5414 10472 5466
rect 10524 5414 10536 5466
rect 10588 5414 10600 5466
rect 10652 5414 10664 5466
rect 10716 5414 10728 5466
rect 10780 5414 19994 5466
rect 20046 5414 20058 5466
rect 20110 5414 20122 5466
rect 20174 5414 20186 5466
rect 20238 5414 20250 5466
rect 20302 5414 29516 5466
rect 29568 5414 29580 5466
rect 29632 5414 29644 5466
rect 29696 5414 29708 5466
rect 29760 5414 29772 5466
rect 29824 5414 39038 5466
rect 39090 5414 39102 5466
rect 39154 5414 39166 5466
rect 39218 5414 39230 5466
rect 39282 5414 39294 5466
rect 39346 5414 39352 5466
rect 1104 5392 39352 5414
rect 1762 5312 1768 5364
rect 1820 5312 1826 5364
rect 6086 5312 6092 5364
rect 6144 5352 6150 5364
rect 8297 5355 8355 5361
rect 6144 5324 8156 5352
rect 6144 5312 6150 5324
rect 2038 5244 2044 5296
rect 2096 5284 2102 5296
rect 2096 5256 3082 5284
rect 2096 5244 2102 5256
rect 4338 5244 4344 5296
rect 4396 5244 4402 5296
rect 5994 5244 6000 5296
rect 6052 5244 6058 5296
rect 7282 5244 7288 5296
rect 7340 5244 7346 5296
rect 8128 5284 8156 5324
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 9398 5352 9404 5364
rect 8343 5324 9404 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 9398 5312 9404 5324
rect 9456 5352 9462 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 9456 5324 9689 5352
rect 9456 5312 9462 5324
rect 9677 5321 9689 5324
rect 9723 5321 9735 5355
rect 9677 5315 9735 5321
rect 10413 5355 10471 5361
rect 10413 5321 10425 5355
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 10428 5284 10456 5315
rect 10962 5312 10968 5364
rect 11020 5352 11026 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 11020 5324 13461 5352
rect 11020 5312 11026 5324
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13449 5315 13507 5321
rect 14001 5355 14059 5361
rect 14001 5321 14013 5355
rect 14047 5352 14059 5355
rect 15010 5352 15016 5364
rect 14047 5324 15016 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 15470 5352 15476 5364
rect 15212 5324 15476 5352
rect 8128 5256 10456 5284
rect 11054 5244 11060 5296
rect 11112 5284 11118 5296
rect 11882 5284 11888 5296
rect 11112 5256 11888 5284
rect 11112 5244 11118 5256
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 13262 5284 13268 5296
rect 13202 5256 13268 5284
rect 13262 5244 13268 5256
rect 13320 5244 13326 5296
rect 13354 5244 13360 5296
rect 13412 5284 13418 5296
rect 15212 5284 15240 5324
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 15654 5312 15660 5364
rect 15712 5352 15718 5364
rect 17862 5352 17868 5364
rect 15712 5324 17868 5352
rect 15712 5312 15718 5324
rect 13412 5256 15240 5284
rect 13412 5244 13418 5256
rect 15286 5244 15292 5296
rect 15344 5244 15350 5296
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 992 5188 1593 5216
rect 992 5176 998 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 5258 5176 5264 5228
rect 5316 5176 5322 5228
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 8996 5188 9536 5216
rect 8996 5176 9002 5188
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5117 2375 5151
rect 2317 5111 2375 5117
rect 1578 5040 1584 5092
rect 1636 5080 1642 5092
rect 2332 5080 2360 5111
rect 2590 5108 2596 5160
rect 2648 5108 2654 5160
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5117 5687 5151
rect 5629 5111 5687 5117
rect 1636 5052 2360 5080
rect 1636 5040 1642 5052
rect 3878 5040 3884 5092
rect 3936 5080 3942 5092
rect 5537 5083 5595 5089
rect 5537 5080 5549 5083
rect 3936 5052 5549 5080
rect 3936 5040 3942 5052
rect 5537 5049 5549 5052
rect 5583 5049 5595 5083
rect 5644 5080 5672 5111
rect 6546 5108 6552 5160
rect 6604 5108 6610 5160
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 9508 5148 9536 5188
rect 9582 5176 9588 5228
rect 9640 5176 9646 5228
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 9692 5188 10793 5216
rect 9692 5148 9720 5188
rect 10781 5185 10793 5188
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5216 13967 5219
rect 14090 5216 14096 5228
rect 13955 5188 14096 5216
rect 13955 5185 13967 5188
rect 13909 5179 13967 5185
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 16868 5225 16896 5324
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18012 5324 20668 5352
rect 18012 5312 18018 5324
rect 17126 5244 17132 5296
rect 17184 5244 17190 5296
rect 17586 5244 17592 5296
rect 17644 5244 17650 5296
rect 18690 5244 18696 5296
rect 18748 5284 18754 5296
rect 18748 5256 19826 5284
rect 18748 5244 18754 5256
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 6871 5120 9260 5148
rect 9508 5120 9720 5148
rect 9769 5151 9827 5157
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 9232 5089 9260 5120
rect 9769 5117 9781 5151
rect 9815 5117 9827 5151
rect 9769 5111 9827 5117
rect 9217 5083 9275 5089
rect 5644 5052 6684 5080
rect 5537 5043 5595 5049
rect 2406 4972 2412 5024
rect 2464 5012 2470 5024
rect 5399 5015 5457 5021
rect 5399 5012 5411 5015
rect 2464 4984 5411 5012
rect 2464 4972 2470 4984
rect 5399 4981 5411 4984
rect 5445 4981 5457 5015
rect 6656 5012 6684 5052
rect 9217 5049 9229 5083
rect 9263 5049 9275 5083
rect 9784 5080 9812 5111
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10192 5120 10885 5148
rect 10192 5108 10198 5120
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 11057 5151 11115 5157
rect 11057 5117 11069 5151
rect 11103 5117 11115 5151
rect 11057 5111 11115 5117
rect 9217 5043 9275 5049
rect 9600 5052 9812 5080
rect 6914 5012 6920 5024
rect 6656 4984 6920 5012
rect 5399 4975 5457 4981
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8202 5012 8208 5024
rect 7984 4984 8208 5012
rect 7984 4972 7990 4984
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 9490 5012 9496 5024
rect 9088 4984 9496 5012
rect 9088 4972 9094 4984
rect 9490 4972 9496 4984
rect 9548 5012 9554 5024
rect 9600 5012 9628 5052
rect 9548 4984 9628 5012
rect 11072 5012 11100 5111
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 11388 5120 11713 5148
rect 11388 5108 11394 5120
rect 11701 5117 11713 5120
rect 11747 5117 11759 5151
rect 11701 5111 11759 5117
rect 11974 5108 11980 5160
rect 12032 5108 12038 5160
rect 14553 5151 14611 5157
rect 14553 5117 14565 5151
rect 14599 5148 14611 5151
rect 14599 5120 14688 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 13906 5012 13912 5024
rect 11072 4984 13912 5012
rect 9548 4972 9554 4984
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14660 5012 14688 5120
rect 14826 5108 14832 5160
rect 14884 5108 14890 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 18601 5151 18659 5157
rect 18601 5148 18613 5151
rect 15436 5120 18613 5148
rect 15436 5108 15442 5120
rect 18601 5117 18613 5120
rect 18647 5117 18659 5151
rect 18601 5111 18659 5117
rect 19058 5108 19064 5160
rect 19116 5108 19122 5160
rect 19337 5151 19395 5157
rect 19337 5148 19349 5151
rect 19168 5120 19349 5148
rect 16114 5040 16120 5092
rect 16172 5080 16178 5092
rect 19168 5080 19196 5120
rect 19337 5117 19349 5120
rect 19383 5117 19395 5151
rect 20640 5148 20668 5324
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 20864 5324 27476 5352
rect 20864 5312 20870 5324
rect 21358 5244 21364 5296
rect 21416 5244 21422 5296
rect 21634 5244 21640 5296
rect 21692 5284 21698 5296
rect 22370 5284 22376 5296
rect 21692 5256 22376 5284
rect 21692 5244 21698 5256
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 22557 5287 22615 5293
rect 22557 5253 22569 5287
rect 22603 5284 22615 5287
rect 22603 5256 22876 5284
rect 22603 5253 22615 5256
rect 22557 5247 22615 5253
rect 21266 5176 21272 5228
rect 21324 5176 21330 5228
rect 22462 5176 22468 5228
rect 22520 5216 22526 5228
rect 22649 5219 22707 5225
rect 22649 5216 22661 5219
rect 22520 5188 22661 5216
rect 22520 5176 22526 5188
rect 22649 5185 22661 5188
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20640 5120 20821 5148
rect 19337 5111 19395 5117
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 20809 5111 20867 5117
rect 22278 5108 22284 5160
rect 22336 5148 22342 5160
rect 22741 5151 22799 5157
rect 22741 5148 22753 5151
rect 22336 5120 22753 5148
rect 22336 5108 22342 5120
rect 22741 5117 22753 5120
rect 22787 5117 22799 5151
rect 22848 5148 22876 5256
rect 23014 5244 23020 5296
rect 23072 5284 23078 5296
rect 23753 5287 23811 5293
rect 23753 5284 23765 5287
rect 23072 5256 23765 5284
rect 23072 5244 23078 5256
rect 23753 5253 23765 5256
rect 23799 5253 23811 5287
rect 25130 5284 25136 5296
rect 23753 5247 23811 5253
rect 24872 5256 25136 5284
rect 22922 5176 22928 5228
rect 22980 5216 22986 5228
rect 22980 5188 23980 5216
rect 22980 5176 22986 5188
rect 22848 5120 23520 5148
rect 22741 5111 22799 5117
rect 16172 5052 16988 5080
rect 16172 5040 16178 5052
rect 14918 5012 14924 5024
rect 14660 4984 14924 5012
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 16298 4972 16304 5024
rect 16356 4972 16362 5024
rect 16960 5012 16988 5052
rect 18892 5052 19196 5080
rect 18892 5012 18920 5052
rect 20346 5040 20352 5092
rect 20404 5080 20410 5092
rect 23385 5083 23443 5089
rect 23385 5080 23397 5083
rect 20404 5052 23397 5080
rect 20404 5040 20410 5052
rect 23385 5049 23397 5052
rect 23431 5049 23443 5083
rect 23492 5080 23520 5120
rect 23842 5108 23848 5160
rect 23900 5108 23906 5160
rect 23952 5157 23980 5188
rect 24670 5176 24676 5228
rect 24728 5216 24734 5228
rect 24872 5225 24900 5256
rect 25130 5244 25136 5256
rect 25188 5244 25194 5296
rect 26878 5284 26884 5296
rect 26358 5256 26884 5284
rect 26878 5244 26884 5256
rect 26936 5244 26942 5296
rect 27338 5244 27344 5296
rect 27396 5244 27402 5296
rect 27448 5284 27476 5324
rect 28166 5312 28172 5364
rect 28224 5352 28230 5364
rect 29362 5352 29368 5364
rect 28224 5324 29368 5352
rect 28224 5312 28230 5324
rect 29362 5312 29368 5324
rect 29420 5312 29426 5364
rect 30282 5312 30288 5364
rect 30340 5352 30346 5364
rect 31665 5355 31723 5361
rect 31665 5352 31677 5355
rect 30340 5324 31677 5352
rect 30340 5312 30346 5324
rect 31665 5321 31677 5324
rect 31711 5321 31723 5355
rect 31665 5315 31723 5321
rect 32122 5312 32128 5364
rect 32180 5352 32186 5364
rect 34698 5352 34704 5364
rect 32180 5324 34704 5352
rect 32180 5312 32186 5324
rect 34698 5312 34704 5324
rect 34756 5312 34762 5364
rect 34790 5312 34796 5364
rect 34848 5352 34854 5364
rect 35345 5355 35403 5361
rect 35345 5352 35357 5355
rect 34848 5324 35357 5352
rect 34848 5312 34854 5324
rect 35345 5321 35357 5324
rect 35391 5321 35403 5355
rect 35345 5315 35403 5321
rect 35710 5312 35716 5364
rect 35768 5352 35774 5364
rect 35805 5355 35863 5361
rect 35805 5352 35817 5355
rect 35768 5324 35817 5352
rect 35768 5312 35774 5324
rect 35805 5321 35817 5324
rect 35851 5321 35863 5355
rect 36630 5352 36636 5364
rect 35805 5315 35863 5321
rect 36464 5324 36636 5352
rect 28534 5284 28540 5296
rect 27448 5256 28540 5284
rect 28534 5244 28540 5256
rect 28592 5244 28598 5296
rect 29914 5244 29920 5296
rect 29972 5284 29978 5296
rect 32585 5287 32643 5293
rect 32585 5284 32597 5287
rect 29972 5256 32597 5284
rect 29972 5244 29978 5256
rect 32585 5253 32597 5256
rect 32631 5253 32643 5287
rect 33502 5284 33508 5296
rect 32585 5247 32643 5253
rect 33152 5256 33508 5284
rect 24857 5219 24915 5225
rect 24857 5216 24869 5219
rect 24728 5188 24869 5216
rect 24728 5176 24734 5188
rect 24857 5185 24869 5188
rect 24903 5185 24915 5219
rect 24857 5179 24915 5185
rect 27157 5219 27215 5225
rect 27157 5185 27169 5219
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27433 5219 27491 5225
rect 27433 5185 27445 5219
rect 27479 5185 27491 5219
rect 27433 5179 27491 5185
rect 23937 5151 23995 5157
rect 23937 5117 23949 5151
rect 23983 5117 23995 5151
rect 23937 5111 23995 5117
rect 24026 5108 24032 5160
rect 24084 5148 24090 5160
rect 25133 5151 25191 5157
rect 25133 5148 25145 5151
rect 24084 5120 25145 5148
rect 24084 5108 24090 5120
rect 25133 5117 25145 5120
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 26605 5151 26663 5157
rect 26605 5117 26617 5151
rect 26651 5148 26663 5151
rect 26970 5148 26976 5160
rect 26651 5120 26976 5148
rect 26651 5117 26663 5120
rect 26605 5111 26663 5117
rect 23492 5052 24164 5080
rect 23385 5043 23443 5049
rect 16960 4984 18920 5012
rect 19058 4972 19064 5024
rect 19116 5012 19122 5024
rect 19426 5012 19432 5024
rect 19116 4984 19432 5012
rect 19116 4972 19122 4984
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 22189 5015 22247 5021
rect 22189 4981 22201 5015
rect 22235 5012 22247 5015
rect 24026 5012 24032 5024
rect 22235 4984 24032 5012
rect 22235 4981 22247 4984
rect 22189 4975 22247 4981
rect 24026 4972 24032 4984
rect 24084 4972 24090 5024
rect 24136 5012 24164 5052
rect 26620 5012 26648 5111
rect 26970 5108 26976 5120
rect 27028 5108 27034 5160
rect 27172 5080 27200 5179
rect 27448 5148 27476 5179
rect 27522 5176 27528 5228
rect 27580 5176 27586 5228
rect 28166 5176 28172 5228
rect 28224 5176 28230 5228
rect 28445 5151 28503 5157
rect 27448 5120 28304 5148
rect 28074 5080 28080 5092
rect 27172 5052 28080 5080
rect 28074 5040 28080 5052
rect 28132 5040 28138 5092
rect 24136 4984 26648 5012
rect 27338 4972 27344 5024
rect 27396 5012 27402 5024
rect 27709 5015 27767 5021
rect 27709 5012 27721 5015
rect 27396 4984 27721 5012
rect 27396 4972 27402 4984
rect 27709 4981 27721 4984
rect 27755 4981 27767 5015
rect 28276 5012 28304 5120
rect 28445 5117 28457 5151
rect 28491 5148 28503 5151
rect 29178 5148 29184 5160
rect 28491 5120 29184 5148
rect 28491 5117 28503 5120
rect 28445 5111 28503 5117
rect 29178 5108 29184 5120
rect 29236 5108 29242 5160
rect 29564 5080 29592 5202
rect 30558 5176 30564 5228
rect 30616 5216 30622 5228
rect 30745 5219 30803 5225
rect 30745 5216 30757 5219
rect 30616 5188 30757 5216
rect 30616 5176 30622 5188
rect 30745 5185 30757 5188
rect 30791 5185 30803 5219
rect 30745 5179 30803 5185
rect 30834 5176 30840 5228
rect 30892 5176 30898 5228
rect 31294 5176 31300 5228
rect 31352 5216 31358 5228
rect 31573 5219 31631 5225
rect 31573 5216 31585 5219
rect 31352 5188 31585 5216
rect 31352 5176 31358 5188
rect 31573 5185 31585 5188
rect 31619 5216 31631 5219
rect 32122 5216 32128 5228
rect 31619 5188 32128 5216
rect 31619 5185 31631 5188
rect 31573 5179 31631 5185
rect 32122 5176 32128 5188
rect 32180 5176 32186 5228
rect 32398 5176 32404 5228
rect 32456 5176 32462 5228
rect 33152 5225 33180 5256
rect 33502 5244 33508 5256
rect 33560 5244 33566 5296
rect 36464 5284 36492 5324
rect 36630 5312 36636 5324
rect 36688 5312 36694 5364
rect 36751 5355 36809 5361
rect 36751 5321 36763 5355
rect 36797 5352 36809 5355
rect 36906 5352 36912 5364
rect 36797 5324 36912 5352
rect 36797 5321 36809 5324
rect 36751 5315 36809 5321
rect 36906 5312 36912 5324
rect 36964 5312 36970 5364
rect 37458 5312 37464 5364
rect 37516 5352 37522 5364
rect 37553 5355 37611 5361
rect 37553 5352 37565 5355
rect 37516 5324 37565 5352
rect 37516 5312 37522 5324
rect 37553 5321 37565 5324
rect 37599 5321 37611 5355
rect 37553 5315 37611 5321
rect 35176 5256 36492 5284
rect 36541 5287 36599 5293
rect 33137 5219 33195 5225
rect 33137 5185 33149 5219
rect 33183 5185 33195 5219
rect 35176 5216 35204 5256
rect 36541 5253 36553 5287
rect 36587 5284 36599 5287
rect 37826 5284 37832 5296
rect 36587 5256 37832 5284
rect 36587 5253 36599 5256
rect 36541 5247 36599 5253
rect 37826 5244 37832 5256
rect 37884 5244 37890 5296
rect 34546 5188 35204 5216
rect 33137 5179 33195 5185
rect 35250 5176 35256 5228
rect 35308 5216 35314 5228
rect 35710 5216 35716 5228
rect 35308 5188 35716 5216
rect 35308 5176 35314 5188
rect 35710 5176 35716 5188
rect 35768 5176 35774 5228
rect 35986 5216 35992 5228
rect 35912 5188 35992 5216
rect 30926 5108 30932 5160
rect 30984 5108 30990 5160
rect 33410 5108 33416 5160
rect 33468 5108 33474 5160
rect 33870 5108 33876 5160
rect 33928 5148 33934 5160
rect 35912 5157 35940 5188
rect 35986 5176 35992 5188
rect 36044 5176 36050 5228
rect 37458 5176 37464 5228
rect 37516 5176 37522 5228
rect 38102 5176 38108 5228
rect 38160 5176 38166 5228
rect 34885 5151 34943 5157
rect 34885 5148 34897 5151
rect 33928 5120 34897 5148
rect 33928 5108 33934 5120
rect 34885 5117 34897 5120
rect 34931 5117 34943 5151
rect 34885 5111 34943 5117
rect 35897 5151 35955 5157
rect 35897 5117 35909 5151
rect 35943 5117 35955 5151
rect 38197 5151 38255 5157
rect 38197 5148 38209 5151
rect 35897 5111 35955 5117
rect 36004 5120 38209 5148
rect 33042 5080 33048 5092
rect 29564 5052 33048 5080
rect 33042 5040 33048 5052
rect 33100 5040 33106 5092
rect 36004 5080 36032 5120
rect 38197 5117 38209 5120
rect 38243 5117 38255 5151
rect 38197 5111 38255 5117
rect 34440 5052 36032 5080
rect 29917 5015 29975 5021
rect 29917 5012 29929 5015
rect 28276 4984 29929 5012
rect 27709 4975 27767 4981
rect 29917 4981 29929 4984
rect 29963 5012 29975 5015
rect 30098 5012 30104 5024
rect 29963 4984 30104 5012
rect 29963 4981 29975 4984
rect 29917 4975 29975 4981
rect 30098 4972 30104 4984
rect 30156 4972 30162 5024
rect 30374 4972 30380 5024
rect 30432 4972 30438 5024
rect 31938 4972 31944 5024
rect 31996 5012 32002 5024
rect 34440 5012 34468 5052
rect 36906 5040 36912 5092
rect 36964 5040 36970 5092
rect 31996 4984 34468 5012
rect 31996 4972 32002 4984
rect 34698 4972 34704 5024
rect 34756 5012 34762 5024
rect 35986 5012 35992 5024
rect 34756 4984 35992 5012
rect 34756 4972 34762 4984
rect 35986 4972 35992 4984
rect 36044 4972 36050 5024
rect 36722 4972 36728 5024
rect 36780 4972 36786 5024
rect 1104 4922 39192 4944
rect 1104 4870 5711 4922
rect 5763 4870 5775 4922
rect 5827 4870 5839 4922
rect 5891 4870 5903 4922
rect 5955 4870 5967 4922
rect 6019 4870 15233 4922
rect 15285 4870 15297 4922
rect 15349 4870 15361 4922
rect 15413 4870 15425 4922
rect 15477 4870 15489 4922
rect 15541 4870 24755 4922
rect 24807 4870 24819 4922
rect 24871 4870 24883 4922
rect 24935 4870 24947 4922
rect 24999 4870 25011 4922
rect 25063 4870 34277 4922
rect 34329 4870 34341 4922
rect 34393 4870 34405 4922
rect 34457 4870 34469 4922
rect 34521 4870 34533 4922
rect 34585 4870 39192 4922
rect 1104 4848 39192 4870
rect 4522 4768 4528 4820
rect 4580 4768 4586 4820
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 4985 4811 5043 4817
rect 4985 4808 4997 4811
rect 4948 4780 4997 4808
rect 4948 4768 4954 4780
rect 4985 4777 4997 4780
rect 5031 4777 5043 4811
rect 4985 4771 5043 4777
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 7929 4811 7987 4817
rect 7929 4808 7941 4811
rect 5132 4780 7941 4808
rect 5132 4768 5138 4780
rect 7929 4777 7941 4780
rect 7975 4777 7987 4811
rect 7929 4771 7987 4777
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 9214 4808 9220 4820
rect 8628 4780 9220 4808
rect 8628 4768 8634 4780
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 9585 4811 9643 4817
rect 9585 4777 9597 4811
rect 9631 4808 9643 4811
rect 11054 4808 11060 4820
rect 9631 4780 11060 4808
rect 9631 4777 9643 4780
rect 9585 4771 9643 4777
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 11425 4811 11483 4817
rect 11425 4777 11437 4811
rect 11471 4808 11483 4811
rect 11974 4808 11980 4820
rect 11471 4780 11980 4808
rect 11471 4777 11483 4780
rect 11425 4771 11483 4777
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 17126 4808 17132 4820
rect 12406 4780 17132 4808
rect 6086 4740 6092 4752
rect 4251 4712 6092 4740
rect 1854 4632 1860 4684
rect 1912 4632 1918 4684
rect 3326 4632 3332 4684
rect 3384 4672 3390 4684
rect 4251 4672 4279 4712
rect 6086 4700 6092 4712
rect 6144 4700 6150 4752
rect 8202 4700 8208 4752
rect 8260 4740 8266 4752
rect 10229 4743 10287 4749
rect 8260 4712 10180 4740
rect 8260 4700 8266 4712
rect 3384 4644 4108 4672
rect 3384 4632 3390 4644
rect 1578 4564 1584 4616
rect 1636 4564 1642 4616
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3752 4576 3985 4604
rect 3752 4564 3758 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 2498 4496 2504 4548
rect 2556 4496 2562 4548
rect 4080 4536 4108 4644
rect 4172 4644 4279 4672
rect 4172 4616 4200 4644
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 5445 4675 5503 4681
rect 5445 4672 5457 4675
rect 5224 4644 5457 4672
rect 5224 4632 5230 4644
rect 5445 4641 5457 4644
rect 5491 4641 5503 4675
rect 5445 4635 5503 4641
rect 5534 4632 5540 4684
rect 5592 4632 5598 4684
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4672 6239 4675
rect 6546 4672 6552 4684
rect 6227 4644 6552 4672
rect 6227 4641 6239 4644
rect 6181 4635 6239 4641
rect 6546 4632 6552 4644
rect 6604 4672 6610 4684
rect 6822 4672 6828 4684
rect 6604 4644 6828 4672
rect 6604 4632 6610 4644
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 9766 4672 9772 4684
rect 8527 4644 9772 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 10152 4672 10180 4712
rect 10229 4709 10241 4743
rect 10275 4740 10287 4743
rect 12406 4740 12434 4780
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 17586 4768 17592 4820
rect 17644 4808 17650 4820
rect 21266 4808 21272 4820
rect 17644 4780 21272 4808
rect 17644 4768 17650 4780
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 22002 4768 22008 4820
rect 22060 4808 22066 4820
rect 22060 4780 24072 4808
rect 22060 4768 22066 4780
rect 10275 4712 12434 4740
rect 12805 4743 12863 4749
rect 10275 4709 10287 4712
rect 10229 4703 10287 4709
rect 12805 4709 12817 4743
rect 12851 4740 12863 4743
rect 14182 4740 14188 4752
rect 12851 4712 14188 4740
rect 12851 4709 12863 4712
rect 12805 4703 12863 4709
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 14734 4740 14740 4752
rect 14292 4712 14740 4740
rect 10870 4672 10876 4684
rect 10152 4644 10876 4672
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 11885 4675 11943 4681
rect 11885 4672 11897 4675
rect 11020 4644 11897 4672
rect 11020 4632 11026 4644
rect 11885 4641 11897 4644
rect 11931 4641 11943 4675
rect 11885 4635 11943 4641
rect 12069 4675 12127 4681
rect 12069 4641 12081 4675
rect 12115 4672 12127 4675
rect 12250 4672 12256 4684
rect 12115 4644 12256 4672
rect 12115 4641 12127 4644
rect 12069 4635 12127 4641
rect 12250 4632 12256 4644
rect 12308 4672 12314 4684
rect 12434 4672 12440 4684
rect 12308 4644 12440 4672
rect 12308 4632 12314 4644
rect 12434 4632 12440 4644
rect 12492 4632 12498 4684
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4672 13323 4675
rect 13354 4672 13360 4684
rect 13311 4644 13360 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 13354 4632 13360 4644
rect 13412 4632 13418 4684
rect 13446 4632 13452 4684
rect 13504 4672 13510 4684
rect 14292 4672 14320 4712
rect 14734 4700 14740 4712
rect 14792 4700 14798 4752
rect 16574 4700 16580 4752
rect 16632 4740 16638 4752
rect 18141 4743 18199 4749
rect 18141 4740 18153 4743
rect 16632 4712 18153 4740
rect 16632 4700 16638 4712
rect 18141 4709 18153 4712
rect 18187 4709 18199 4743
rect 20530 4740 20536 4752
rect 18141 4703 18199 4709
rect 18800 4712 20536 4740
rect 13504 4644 14320 4672
rect 13504 4632 13510 4644
rect 14550 4632 14556 4684
rect 14608 4672 14614 4684
rect 14608 4644 14688 4672
rect 14608 4632 14614 4644
rect 4154 4564 4160 4616
rect 4212 4564 4218 4616
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 5902 4604 5908 4616
rect 4387 4576 5908 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 8352 4576 8401 4604
rect 8352 4564 8358 4576
rect 8389 4573 8401 4576
rect 8435 4604 8447 4607
rect 8570 4604 8576 4616
rect 8435 4576 8576 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4573 9091 4607
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 9033 4567 9091 4573
rect 9140 4576 9413 4604
rect 4080 4508 5475 4536
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 5074 4468 5080 4480
rect 4672 4440 5080 4468
rect 4672 4428 4678 4440
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 5353 4471 5411 4477
rect 5353 4468 5365 4471
rect 5224 4440 5365 4468
rect 5224 4428 5230 4440
rect 5353 4437 5365 4440
rect 5399 4437 5411 4471
rect 5447 4468 5475 4508
rect 5718 4496 5724 4548
rect 5776 4536 5782 4548
rect 6457 4539 6515 4545
rect 6457 4536 6469 4539
rect 5776 4508 6469 4536
rect 5776 4496 5782 4508
rect 6457 4505 6469 4508
rect 6503 4505 6515 4539
rect 7742 4536 7748 4548
rect 7682 4508 7748 4536
rect 6457 4499 6515 4505
rect 7742 4496 7748 4508
rect 7800 4496 7806 4548
rect 9048 4536 9076 4567
rect 7852 4508 9076 4536
rect 7852 4468 7880 4508
rect 5447 4440 7880 4468
rect 5353 4431 5411 4437
rect 7926 4428 7932 4480
rect 7984 4468 7990 4480
rect 9140 4468 9168 4576
rect 9401 4573 9413 4576
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9732 4576 9873 4604
rect 9732 4564 9738 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 11146 4604 11152 4616
rect 9861 4567 9919 4573
rect 10612 4576 11152 4604
rect 9214 4496 9220 4548
rect 9272 4496 9278 4548
rect 9309 4539 9367 4545
rect 9309 4505 9321 4539
rect 9355 4536 9367 4539
rect 10612 4536 10640 4576
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 12986 4604 12992 4616
rect 11296 4576 12992 4604
rect 11296 4564 11302 4576
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13964 4576 14289 4604
rect 13964 4564 13970 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 14458 4564 14464 4616
rect 14516 4564 14522 4616
rect 14660 4613 14688 4644
rect 14918 4632 14924 4684
rect 14976 4672 14982 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 14976 4644 15301 4672
rect 14976 4632 14982 4644
rect 15289 4641 15301 4644
rect 15335 4672 15347 4675
rect 15654 4672 15660 4684
rect 15335 4644 15660 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 17037 4675 17095 4681
rect 17037 4641 17049 4675
rect 17083 4672 17095 4675
rect 17678 4672 17684 4684
rect 17083 4644 17684 4672
rect 17083 4641 17095 4644
rect 17037 4635 17095 4641
rect 17678 4632 17684 4644
rect 17736 4632 17742 4684
rect 18322 4632 18328 4684
rect 18380 4672 18386 4684
rect 18800 4681 18828 4712
rect 20530 4700 20536 4712
rect 20588 4700 20594 4752
rect 22186 4700 22192 4752
rect 22244 4740 22250 4752
rect 22922 4740 22928 4752
rect 22244 4712 22928 4740
rect 22244 4700 22250 4712
rect 22922 4700 22928 4712
rect 22980 4700 22986 4752
rect 23934 4740 23940 4752
rect 23308 4712 23940 4740
rect 18601 4675 18659 4681
rect 18601 4672 18613 4675
rect 18380 4644 18613 4672
rect 18380 4632 18386 4644
rect 18601 4641 18613 4644
rect 18647 4641 18659 4675
rect 18601 4635 18659 4641
rect 18785 4675 18843 4681
rect 18785 4641 18797 4675
rect 18831 4641 18843 4675
rect 18785 4635 18843 4641
rect 19886 4632 19892 4684
rect 19944 4632 19950 4684
rect 19978 4632 19984 4684
rect 20036 4632 20042 4684
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 22646 4672 22652 4684
rect 20947 4644 22652 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 22646 4632 22652 4644
rect 22704 4632 22710 4684
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4573 14703 4607
rect 14645 4567 14703 4573
rect 9355 4508 10640 4536
rect 10689 4539 10747 4545
rect 9355 4505 9367 4508
rect 9309 4499 9367 4505
rect 10689 4505 10701 4539
rect 10735 4536 10747 4539
rect 10735 4508 14320 4536
rect 10735 4505 10747 4508
rect 10689 4499 10747 4505
rect 14292 4480 14320 4508
rect 14550 4496 14556 4548
rect 14608 4496 14614 4548
rect 14660 4536 14688 4567
rect 16666 4564 16672 4616
rect 16724 4564 16730 4616
rect 16942 4564 16948 4616
rect 17000 4604 17006 4616
rect 17000 4576 19380 4604
rect 17000 4564 17006 4576
rect 15470 4536 15476 4548
rect 14660 4508 15476 4536
rect 15470 4496 15476 4508
rect 15528 4496 15534 4548
rect 15562 4496 15568 4548
rect 15620 4496 15626 4548
rect 19242 4536 19248 4548
rect 17144 4508 19248 4536
rect 7984 4440 9168 4468
rect 7984 4428 7990 4440
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10597 4471 10655 4477
rect 10597 4468 10609 4471
rect 9732 4440 10609 4468
rect 9732 4428 9738 4440
rect 10597 4437 10609 4440
rect 10643 4437 10655 4471
rect 10597 4431 10655 4437
rect 11793 4471 11851 4477
rect 11793 4437 11805 4471
rect 11839 4468 11851 4471
rect 12158 4468 12164 4480
rect 11839 4440 12164 4468
rect 11839 4437 11851 4440
rect 11793 4431 11851 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 13170 4428 13176 4480
rect 13228 4428 13234 4480
rect 14274 4428 14280 4480
rect 14332 4428 14338 4480
rect 14829 4471 14887 4477
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 17144 4468 17172 4508
rect 19242 4496 19248 4508
rect 19300 4496 19306 4548
rect 19352 4536 19380 4576
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 20622 4604 20628 4616
rect 19484 4576 20628 4604
rect 19484 4564 19490 4576
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 22830 4564 22836 4616
rect 22888 4604 22894 4616
rect 23198 4604 23204 4616
rect 22888 4576 23204 4604
rect 22888 4564 22894 4576
rect 23198 4564 23204 4576
rect 23256 4564 23262 4616
rect 22649 4539 22707 4545
rect 19352 4508 21390 4536
rect 22649 4505 22661 4539
rect 22695 4536 22707 4539
rect 23308 4536 23336 4712
rect 23934 4700 23940 4712
rect 23992 4700 23998 4752
rect 24044 4740 24072 4780
rect 25774 4768 25780 4820
rect 25832 4768 25838 4820
rect 26050 4768 26056 4820
rect 26108 4768 26114 4820
rect 27430 4808 27436 4820
rect 26896 4780 27436 4808
rect 26145 4743 26203 4749
rect 26145 4740 26157 4743
rect 24044 4712 26157 4740
rect 26145 4709 26157 4712
rect 26191 4709 26203 4743
rect 26145 4703 26203 4709
rect 23382 4632 23388 4684
rect 23440 4672 23446 4684
rect 26237 4675 26295 4681
rect 26237 4672 26249 4675
rect 23440 4644 26249 4672
rect 23440 4632 23446 4644
rect 26237 4641 26249 4644
rect 26283 4641 26295 4675
rect 26237 4635 26295 4641
rect 23566 4564 23572 4616
rect 23624 4564 23630 4616
rect 24394 4564 24400 4616
rect 24452 4604 24458 4616
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 24452 4576 24685 4604
rect 24452 4564 24458 4576
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 26326 4564 26332 4616
rect 26384 4564 26390 4616
rect 26513 4607 26571 4613
rect 26513 4573 26525 4607
rect 26559 4604 26571 4607
rect 26896 4604 26924 4780
rect 27430 4768 27436 4780
rect 27488 4768 27494 4820
rect 28994 4768 29000 4820
rect 29052 4808 29058 4820
rect 30098 4808 30104 4820
rect 29052 4780 30104 4808
rect 29052 4768 29058 4780
rect 30098 4768 30104 4780
rect 30156 4808 30162 4820
rect 33781 4811 33839 4817
rect 33781 4808 33793 4811
rect 30156 4780 33793 4808
rect 30156 4768 30162 4780
rect 33781 4777 33793 4780
rect 33827 4777 33839 4811
rect 33781 4771 33839 4777
rect 34422 4768 34428 4820
rect 34480 4808 34486 4820
rect 36170 4808 36176 4820
rect 34480 4780 36176 4808
rect 34480 4768 34486 4780
rect 36170 4768 36176 4780
rect 36228 4768 36234 4820
rect 36538 4768 36544 4820
rect 36596 4808 36602 4820
rect 36633 4811 36691 4817
rect 36633 4808 36645 4811
rect 36596 4780 36645 4808
rect 36596 4768 36602 4780
rect 36633 4777 36645 4780
rect 36679 4777 36691 4811
rect 36633 4771 36691 4777
rect 37182 4768 37188 4820
rect 37240 4808 37246 4820
rect 38565 4811 38623 4817
rect 38565 4808 38577 4811
rect 37240 4780 38577 4808
rect 37240 4768 37246 4780
rect 38565 4777 38577 4780
rect 38611 4777 38623 4811
rect 38565 4771 38623 4777
rect 26973 4743 27031 4749
rect 26973 4709 26985 4743
rect 27019 4740 27031 4743
rect 27019 4712 29316 4740
rect 27019 4709 27031 4712
rect 26973 4703 27031 4709
rect 27246 4632 27252 4684
rect 27304 4672 27310 4684
rect 27525 4675 27583 4681
rect 27525 4672 27537 4675
rect 27304 4644 27537 4672
rect 27304 4632 27310 4644
rect 27525 4641 27537 4644
rect 27571 4641 27583 4675
rect 28994 4672 29000 4684
rect 27525 4635 27583 4641
rect 27632 4644 29000 4672
rect 26559 4576 26924 4604
rect 27433 4607 27491 4613
rect 26559 4573 26571 4576
rect 26513 4567 26571 4573
rect 27433 4573 27445 4607
rect 27479 4604 27491 4607
rect 27632 4604 27660 4644
rect 28994 4632 29000 4644
rect 29052 4632 29058 4684
rect 27479 4576 27660 4604
rect 27479 4573 27491 4576
rect 27433 4567 27491 4573
rect 28166 4564 28172 4616
rect 28224 4564 28230 4616
rect 28350 4564 28356 4616
rect 28408 4564 28414 4616
rect 28534 4564 28540 4616
rect 28592 4564 28598 4616
rect 22695 4508 23336 4536
rect 22695 4505 22707 4508
rect 22649 4499 22707 4505
rect 23474 4496 23480 4548
rect 23532 4536 23538 4548
rect 23842 4536 23848 4548
rect 23532 4508 23848 4536
rect 23532 4496 23538 4508
rect 23842 4496 23848 4508
rect 23900 4536 23906 4548
rect 24762 4536 24768 4548
rect 23900 4508 24768 4536
rect 23900 4496 23906 4508
rect 24762 4496 24768 4508
rect 24820 4496 24826 4548
rect 25225 4539 25283 4545
rect 25225 4505 25237 4539
rect 25271 4536 25283 4539
rect 25774 4536 25780 4548
rect 25271 4508 25780 4536
rect 25271 4505 25283 4508
rect 25225 4499 25283 4505
rect 14875 4440 17172 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 18506 4428 18512 4480
rect 18564 4428 18570 4480
rect 19429 4471 19487 4477
rect 19429 4437 19441 4471
rect 19475 4468 19487 4471
rect 19610 4468 19616 4480
rect 19475 4440 19616 4468
rect 19475 4437 19487 4440
rect 19429 4431 19487 4437
rect 19610 4428 19616 4440
rect 19668 4428 19674 4480
rect 19797 4471 19855 4477
rect 19797 4437 19809 4471
rect 19843 4468 19855 4471
rect 20254 4468 20260 4480
rect 19843 4440 20260 4468
rect 19843 4437 19855 4440
rect 19797 4431 19855 4437
rect 20254 4428 20260 4440
rect 20312 4428 20318 4480
rect 21266 4428 21272 4480
rect 21324 4468 21330 4480
rect 25240 4468 25268 4499
rect 25774 4496 25780 4508
rect 25832 4496 25838 4548
rect 26234 4496 26240 4548
rect 26292 4536 26298 4548
rect 27341 4539 27399 4545
rect 27341 4536 27353 4539
rect 26292 4508 27353 4536
rect 26292 4496 26298 4508
rect 27341 4505 27353 4508
rect 27387 4536 27399 4539
rect 28258 4536 28264 4548
rect 27387 4508 28264 4536
rect 27387 4505 27399 4508
rect 27341 4499 27399 4505
rect 28258 4496 28264 4508
rect 28316 4496 28322 4548
rect 28442 4496 28448 4548
rect 28500 4496 28506 4548
rect 21324 4440 25268 4468
rect 21324 4428 21330 4440
rect 27522 4428 27528 4480
rect 27580 4468 27586 4480
rect 28721 4471 28779 4477
rect 28721 4468 28733 4471
rect 27580 4440 28733 4468
rect 27580 4428 27586 4440
rect 28721 4437 28733 4440
rect 28767 4437 28779 4471
rect 29288 4468 29316 4712
rect 31018 4700 31024 4752
rect 31076 4740 31082 4752
rect 31481 4743 31539 4749
rect 31481 4740 31493 4743
rect 31076 4712 31493 4740
rect 31076 4700 31082 4712
rect 31481 4709 31493 4712
rect 31527 4709 31539 4743
rect 37277 4743 37335 4749
rect 37277 4740 37289 4743
rect 31481 4703 31539 4709
rect 33336 4712 37289 4740
rect 30006 4632 30012 4684
rect 30064 4632 30070 4684
rect 32030 4632 32036 4684
rect 32088 4632 32094 4684
rect 33042 4632 33048 4684
rect 33100 4672 33106 4684
rect 33336 4672 33364 4712
rect 37277 4709 37289 4712
rect 37323 4709 37335 4743
rect 37277 4703 37335 4709
rect 37921 4675 37979 4681
rect 37921 4672 37933 4675
rect 33100 4644 33364 4672
rect 33428 4644 37933 4672
rect 33100 4632 33106 4644
rect 29362 4564 29368 4616
rect 29420 4604 29426 4616
rect 29733 4607 29791 4613
rect 29733 4604 29745 4607
rect 29420 4576 29745 4604
rect 29420 4564 29426 4576
rect 29733 4573 29745 4576
rect 29779 4573 29791 4607
rect 31938 4604 31944 4616
rect 31142 4576 31944 4604
rect 29733 4567 29791 4573
rect 31938 4564 31944 4576
rect 31996 4564 32002 4616
rect 33428 4590 33456 4644
rect 37921 4641 37933 4644
rect 37967 4641 37979 4675
rect 37921 4635 37979 4641
rect 35066 4564 35072 4616
rect 35124 4604 35130 4616
rect 35437 4607 35495 4613
rect 35437 4604 35449 4607
rect 35124 4576 35449 4604
rect 35124 4564 35130 4576
rect 35437 4573 35449 4576
rect 35483 4573 35495 4607
rect 35437 4567 35495 4573
rect 36170 4564 36176 4616
rect 36228 4604 36234 4616
rect 36541 4607 36599 4613
rect 36541 4604 36553 4607
rect 36228 4576 36553 4604
rect 36228 4564 36234 4576
rect 36541 4573 36553 4576
rect 36587 4573 36599 4607
rect 36541 4567 36599 4573
rect 30006 4496 30012 4548
rect 30064 4536 30070 4548
rect 30282 4536 30288 4548
rect 30064 4508 30288 4536
rect 30064 4496 30070 4508
rect 30282 4496 30288 4508
rect 30340 4496 30346 4548
rect 32309 4539 32367 4545
rect 32309 4536 32321 4539
rect 31312 4508 32321 4536
rect 31312 4468 31340 4508
rect 32309 4505 32321 4508
rect 32355 4505 32367 4539
rect 32309 4499 32367 4505
rect 33778 4496 33784 4548
rect 33836 4536 33842 4548
rect 35805 4539 35863 4545
rect 35805 4536 35817 4539
rect 33836 4508 35817 4536
rect 33836 4496 33842 4508
rect 35805 4505 35817 4508
rect 35851 4505 35863 4539
rect 36556 4536 36584 4567
rect 37182 4564 37188 4616
rect 37240 4564 37246 4616
rect 37550 4604 37556 4616
rect 37292 4576 37556 4604
rect 37090 4536 37096 4548
rect 36556 4508 37096 4536
rect 35805 4499 35863 4505
rect 37090 4496 37096 4508
rect 37148 4536 37154 4548
rect 37292 4536 37320 4576
rect 37550 4564 37556 4576
rect 37608 4604 37614 4616
rect 37829 4607 37887 4613
rect 37829 4604 37841 4607
rect 37608 4576 37841 4604
rect 37608 4564 37614 4576
rect 37829 4573 37841 4576
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 38473 4607 38531 4613
rect 38473 4573 38485 4607
rect 38519 4573 38531 4607
rect 38473 4567 38531 4573
rect 37148 4508 37320 4536
rect 37148 4496 37154 4508
rect 37458 4496 37464 4548
rect 37516 4536 37522 4548
rect 38378 4536 38384 4548
rect 37516 4508 38384 4536
rect 37516 4496 37522 4508
rect 38378 4496 38384 4508
rect 38436 4536 38442 4548
rect 38488 4536 38516 4567
rect 38436 4508 38516 4536
rect 38436 4496 38442 4508
rect 29288 4440 31340 4468
rect 28721 4431 28779 4437
rect 32122 4428 32128 4480
rect 32180 4468 32186 4480
rect 34422 4468 34428 4480
rect 32180 4440 34428 4468
rect 32180 4428 32186 4440
rect 34422 4428 34428 4440
rect 34480 4428 34486 4480
rect 34790 4428 34796 4480
rect 34848 4468 34854 4480
rect 38286 4468 38292 4480
rect 34848 4440 38292 4468
rect 34848 4428 34854 4440
rect 38286 4428 38292 4440
rect 38344 4428 38350 4480
rect 1104 4378 39352 4400
rect 1104 4326 10472 4378
rect 10524 4326 10536 4378
rect 10588 4326 10600 4378
rect 10652 4326 10664 4378
rect 10716 4326 10728 4378
rect 10780 4326 19994 4378
rect 20046 4326 20058 4378
rect 20110 4326 20122 4378
rect 20174 4326 20186 4378
rect 20238 4326 20250 4378
rect 20302 4326 29516 4378
rect 29568 4326 29580 4378
rect 29632 4326 29644 4378
rect 29696 4326 29708 4378
rect 29760 4326 29772 4378
rect 29824 4326 39038 4378
rect 39090 4326 39102 4378
rect 39154 4326 39166 4378
rect 39218 4326 39230 4378
rect 39282 4326 39294 4378
rect 39346 4326 39352 4378
rect 1104 4304 39352 4326
rect 5442 4264 5448 4276
rect 2746 4236 5448 4264
rect 1673 4199 1731 4205
rect 1673 4165 1685 4199
rect 1719 4196 1731 4199
rect 2746 4196 2774 4236
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 5629 4267 5687 4273
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 8021 4267 8079 4273
rect 8021 4264 8033 4267
rect 5675 4236 8033 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 8021 4233 8033 4236
rect 8067 4264 8079 4267
rect 8478 4264 8484 4276
rect 8067 4236 8484 4264
rect 8067 4233 8079 4236
rect 8021 4227 8079 4233
rect 1719 4168 2774 4196
rect 1719 4165 1731 4168
rect 1673 4159 1731 4165
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 3016 4168 3542 4196
rect 3016 4156 3022 4168
rect 5166 4156 5172 4208
rect 5224 4196 5230 4208
rect 5644 4196 5672 4227
rect 8478 4224 8484 4236
rect 8536 4224 8542 4276
rect 9217 4267 9275 4273
rect 9217 4233 9229 4267
rect 9263 4264 9275 4267
rect 13354 4264 13360 4276
rect 9263 4236 13360 4264
rect 9263 4233 9275 4236
rect 9217 4227 9275 4233
rect 13354 4224 13360 4236
rect 13412 4264 13418 4276
rect 13906 4264 13912 4276
rect 13412 4236 13912 4264
rect 13412 4224 13418 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14056 4236 17724 4264
rect 14056 4224 14062 4236
rect 5224 4168 5672 4196
rect 5224 4156 5230 4168
rect 5902 4156 5908 4208
rect 5960 4196 5966 4208
rect 5960 4168 7052 4196
rect 5960 4156 5966 4168
rect 5626 4128 5632 4140
rect 4448 4100 5632 4128
rect 1578 4020 1584 4072
rect 1636 4060 1642 4072
rect 2777 4063 2835 4069
rect 2777 4060 2789 4063
rect 1636 4032 2789 4060
rect 1636 4020 1642 4032
rect 2777 4029 2789 4032
rect 2823 4029 2835 4063
rect 2777 4023 2835 4029
rect 3050 4020 3056 4072
rect 3108 4020 3114 4072
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 4448 4060 4476 4100
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 6638 4088 6644 4140
rect 6696 4088 6702 4140
rect 7024 4137 7052 4168
rect 7282 4156 7288 4208
rect 7340 4196 7346 4208
rect 8202 4196 8208 4208
rect 7340 4168 8208 4196
rect 7340 4156 7346 4168
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 10318 4156 10324 4208
rect 10376 4196 10382 4208
rect 10597 4199 10655 4205
rect 10597 4196 10609 4199
rect 10376 4168 10609 4196
rect 10376 4156 10382 4168
rect 10597 4165 10609 4168
rect 10643 4165 10655 4199
rect 10597 4159 10655 4165
rect 10686 4156 10692 4208
rect 10744 4196 10750 4208
rect 13446 4196 13452 4208
rect 10744 4168 13452 4196
rect 10744 4156 10750 4168
rect 13446 4156 13452 4168
rect 13504 4156 13510 4208
rect 14826 4196 14832 4208
rect 14292 4168 14832 4196
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4128 7067 4131
rect 7098 4128 7104 4140
rect 7055 4100 7104 4128
rect 7055 4097 7067 4100
rect 7009 4091 7067 4097
rect 3476 4032 4476 4060
rect 3476 4020 3482 4032
rect 4522 4020 4528 4072
rect 4580 4020 4586 4072
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 5810 4060 5816 4072
rect 5767 4032 5816 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 5902 4020 5908 4072
rect 5960 4020 5966 4072
rect 6546 4020 6552 4072
rect 6604 4060 6610 4072
rect 6840 4060 6868 4091
rect 6604 4032 6868 4060
rect 6932 4060 6960 4091
rect 7098 4088 7104 4100
rect 7156 4128 7162 4140
rect 7926 4128 7932 4140
rect 7156 4100 7932 4128
rect 7156 4088 7162 4100
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 8110 4060 8116 4072
rect 6932 4032 7052 4060
rect 6604 4020 6610 4032
rect 7024 4004 7052 4032
rect 7116 4032 8116 4060
rect 4338 3952 4344 4004
rect 4396 3992 4402 4004
rect 4396 3964 6960 3992
rect 4396 3952 4402 3964
rect 1762 3884 1768 3936
rect 1820 3884 1826 3936
rect 5261 3927 5319 3933
rect 5261 3893 5273 3927
rect 5307 3924 5319 3927
rect 5350 3924 5356 3936
rect 5307 3896 5356 3924
rect 5307 3893 5319 3896
rect 5261 3887 5319 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 6730 3924 6736 3936
rect 5684 3896 6736 3924
rect 5684 3884 5690 3896
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 6932 3924 6960 3964
rect 7006 3952 7012 4004
rect 7064 3952 7070 4004
rect 7116 3924 7144 4032
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8220 4069 8248 4156
rect 14292 4140 14320 4168
rect 14826 4156 14832 4168
rect 14884 4156 14890 4208
rect 15194 4156 15200 4208
rect 15252 4156 15258 4208
rect 17586 4196 17592 4208
rect 15856 4168 17592 4196
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4128 9367 4131
rect 10226 4128 10232 4140
rect 9355 4100 10232 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 11701 4131 11759 4137
rect 10428 4100 10824 4128
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 9674 4060 9680 4072
rect 9539 4032 9680 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 9674 4020 9680 4032
rect 9732 4060 9738 4072
rect 10134 4060 10140 4072
rect 9732 4032 10140 4060
rect 9732 4020 9738 4032
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 10428 4060 10456 4100
rect 10244 4032 10456 4060
rect 10597 4063 10655 4069
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 10244 3992 10272 4032
rect 10597 4029 10609 4063
rect 10643 4029 10655 4063
rect 10796 4060 10824 4100
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 12066 4128 12072 4140
rect 11747 4100 12072 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12342 4088 12348 4140
rect 12400 4088 12406 4140
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12544 4060 12572 4091
rect 12894 4088 12900 4140
rect 12952 4088 12958 4140
rect 13078 4088 13084 4140
rect 13136 4088 13142 4140
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 10796 4032 12572 4060
rect 10597 4023 10655 4029
rect 7239 3964 10272 3992
rect 10612 3992 10640 4023
rect 12986 4020 12992 4072
rect 13044 4060 13050 4072
rect 13280 4060 13308 4091
rect 14274 4088 14280 4140
rect 14332 4088 14338 4140
rect 13044 4032 13308 4060
rect 13044 4020 13050 4032
rect 14182 4020 14188 4072
rect 14240 4060 14246 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 14240 4032 14565 4060
rect 14240 4020 14246 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 15562 4060 15568 4072
rect 14700 4032 15568 4060
rect 14700 4020 14706 4032
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 15856 4060 15884 4168
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 17696 4196 17724 4236
rect 20438 4224 20444 4276
rect 20496 4264 20502 4276
rect 20496 4236 22094 4264
rect 20496 4224 20502 4236
rect 17696 4168 18722 4196
rect 19518 4156 19524 4208
rect 19576 4196 19582 4208
rect 19576 4168 20760 4196
rect 19576 4156 19582 4168
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 15672 4032 15884 4060
rect 16960 4060 16988 4091
rect 17034 4088 17040 4140
rect 17092 4128 17098 4140
rect 17129 4131 17187 4137
rect 17129 4128 17141 4131
rect 17092 4100 17141 4128
rect 17092 4088 17098 4100
rect 17129 4097 17141 4100
rect 17175 4097 17187 4131
rect 17129 4091 17187 4097
rect 17218 4088 17224 4140
rect 17276 4088 17282 4140
rect 17310 4088 17316 4140
rect 17368 4088 17374 4140
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 17957 4131 18015 4137
rect 17957 4128 17969 4131
rect 17920 4100 17969 4128
rect 17920 4088 17926 4100
rect 17957 4097 17969 4100
rect 18003 4097 18015 4131
rect 20732 4128 20760 4168
rect 20990 4156 20996 4208
rect 21048 4196 21054 4208
rect 21085 4199 21143 4205
rect 21085 4196 21097 4199
rect 21048 4168 21097 4196
rect 21048 4156 21054 4168
rect 21085 4165 21097 4168
rect 21131 4165 21143 4199
rect 22066 4196 22094 4236
rect 22278 4224 22284 4276
rect 22336 4264 22342 4276
rect 22922 4264 22928 4276
rect 22336 4236 22928 4264
rect 22336 4224 22342 4236
rect 22922 4224 22928 4236
rect 22980 4224 22986 4276
rect 24029 4267 24087 4273
rect 24029 4233 24041 4267
rect 24075 4233 24087 4267
rect 24029 4227 24087 4233
rect 22066 4168 23046 4196
rect 21085 4159 21143 4165
rect 24044 4140 24072 4227
rect 24486 4224 24492 4276
rect 24544 4264 24550 4276
rect 24949 4267 25007 4273
rect 24949 4264 24961 4267
rect 24544 4236 24961 4264
rect 24544 4224 24550 4236
rect 24949 4233 24961 4236
rect 24995 4233 25007 4267
rect 24949 4227 25007 4233
rect 26053 4267 26111 4273
rect 26053 4233 26065 4267
rect 26099 4264 26111 4267
rect 26234 4264 26240 4276
rect 26099 4236 26240 4264
rect 26099 4233 26111 4236
rect 26053 4227 26111 4233
rect 26234 4224 26240 4236
rect 26292 4224 26298 4276
rect 28166 4224 28172 4276
rect 28224 4264 28230 4276
rect 31938 4264 31944 4276
rect 28224 4236 31944 4264
rect 28224 4224 28230 4236
rect 31938 4224 31944 4236
rect 31996 4224 32002 4276
rect 35158 4264 35164 4276
rect 32968 4236 35164 4264
rect 24780 4168 24992 4196
rect 21177 4131 21235 4137
rect 21177 4128 21189 4131
rect 20732 4100 21189 4128
rect 17957 4091 18015 4097
rect 21177 4097 21189 4100
rect 21223 4128 21235 4131
rect 21634 4128 21640 4140
rect 21223 4100 21640 4128
rect 21223 4097 21235 4100
rect 21177 4091 21235 4097
rect 21634 4088 21640 4100
rect 21692 4088 21698 4140
rect 24026 4088 24032 4140
rect 24084 4128 24090 4140
rect 24780 4128 24808 4168
rect 24084 4100 24808 4128
rect 24084 4088 24090 4100
rect 24854 4088 24860 4140
rect 24912 4088 24918 4140
rect 24964 4128 24992 4168
rect 25976 4168 26188 4196
rect 25976 4128 26004 4168
rect 24964 4100 26004 4128
rect 26160 4128 26188 4168
rect 26602 4156 26608 4208
rect 26660 4196 26666 4208
rect 26660 4168 27384 4196
rect 26660 4156 26666 4168
rect 27356 4137 27384 4168
rect 28074 4156 28080 4208
rect 28132 4196 28138 4208
rect 30006 4196 30012 4208
rect 28132 4168 28488 4196
rect 28132 4156 28138 4168
rect 28460 4137 28488 4168
rect 28828 4168 30012 4196
rect 27341 4131 27399 4137
rect 26160 4100 27292 4128
rect 17770 4060 17776 4072
rect 16960 4032 17776 4060
rect 12802 3992 12808 4004
rect 10612 3964 11928 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 6932 3896 7144 3924
rect 7650 3884 7656 3936
rect 7708 3884 7714 3936
rect 8846 3884 8852 3936
rect 8904 3884 8910 3936
rect 10134 3884 10140 3936
rect 10192 3884 10198 3936
rect 11790 3884 11796 3936
rect 11848 3884 11854 3936
rect 11900 3924 11928 3964
rect 12636 3964 12808 3992
rect 12636 3924 12664 3964
rect 12802 3952 12808 3964
rect 12860 3992 12866 4004
rect 13906 3992 13912 4004
rect 12860 3964 13912 3992
rect 12860 3952 12866 3964
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 11900 3896 12664 3924
rect 13630 3884 13636 3936
rect 13688 3924 13694 3936
rect 13725 3927 13783 3933
rect 13725 3924 13737 3927
rect 13688 3896 13737 3924
rect 13688 3884 13694 3896
rect 13725 3893 13737 3896
rect 13771 3893 13783 3927
rect 13725 3887 13783 3893
rect 14090 3884 14096 3936
rect 14148 3924 14154 3936
rect 15672 3924 15700 4032
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 17126 3952 17132 4004
rect 17184 3992 17190 4004
rect 17880 3992 17908 4088
rect 18233 4063 18291 4069
rect 18233 4029 18245 4063
rect 18279 4060 18291 4063
rect 20346 4060 20352 4072
rect 18279 4032 20352 4060
rect 18279 4029 18291 4032
rect 18233 4023 18291 4029
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 21358 4020 21364 4072
rect 21416 4020 21422 4072
rect 22281 4063 22339 4069
rect 22281 4029 22293 4063
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 17184 3964 17908 3992
rect 17184 3952 17190 3964
rect 19334 3952 19340 4004
rect 19392 3992 19398 4004
rect 19705 3995 19763 4001
rect 19705 3992 19717 3995
rect 19392 3964 19717 3992
rect 19392 3952 19398 3964
rect 19705 3961 19717 3964
rect 19751 3961 19763 3995
rect 19705 3955 19763 3961
rect 20622 3952 20628 4004
rect 20680 3992 20686 4004
rect 22296 3992 22324 4023
rect 22554 4020 22560 4072
rect 22612 4020 22618 4072
rect 22646 4020 22652 4072
rect 22704 4060 22710 4072
rect 22704 4032 24900 4060
rect 22704 4020 22710 4032
rect 24670 3992 24676 4004
rect 20680 3964 22324 3992
rect 20680 3952 20686 3964
rect 14148 3896 15700 3924
rect 14148 3884 14154 3896
rect 15746 3884 15752 3936
rect 15804 3924 15810 3936
rect 17310 3924 17316 3936
rect 15804 3896 17316 3924
rect 15804 3884 15810 3896
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 17497 3927 17555 3933
rect 17497 3893 17509 3927
rect 17543 3924 17555 3927
rect 19518 3924 19524 3936
rect 17543 3896 19524 3924
rect 17543 3893 17555 3896
rect 17497 3887 17555 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 20717 3927 20775 3933
rect 20717 3893 20729 3927
rect 20763 3924 20775 3927
rect 22186 3924 22192 3936
rect 20763 3896 22192 3924
rect 20763 3893 20775 3896
rect 20717 3887 20775 3893
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 22296 3924 22324 3964
rect 23584 3964 24676 3992
rect 23584 3924 23612 3964
rect 24670 3952 24676 3964
rect 24728 3952 24734 4004
rect 24872 3992 24900 4032
rect 25130 4020 25136 4072
rect 25188 4020 25194 4072
rect 26145 4063 26203 4069
rect 26145 4029 26157 4063
rect 26191 4029 26203 4063
rect 26145 4023 26203 4029
rect 26160 3992 26188 4023
rect 26234 4020 26240 4072
rect 26292 4020 26298 4072
rect 27157 4063 27215 4069
rect 27157 4029 27169 4063
rect 27203 4029 27215 4063
rect 27264 4060 27292 4100
rect 27341 4097 27353 4131
rect 27387 4097 27399 4131
rect 27341 4091 27399 4097
rect 28353 4131 28411 4137
rect 28353 4097 28365 4131
rect 28399 4097 28411 4131
rect 28353 4091 28411 4097
rect 28445 4131 28503 4137
rect 28445 4097 28457 4131
rect 28491 4128 28503 4131
rect 28718 4128 28724 4140
rect 28491 4100 28724 4128
rect 28491 4097 28503 4100
rect 28445 4091 28503 4097
rect 27264 4032 28120 4060
rect 27157 4023 27215 4029
rect 27172 3992 27200 4023
rect 24872 3964 27200 3992
rect 22296 3896 23612 3924
rect 24486 3884 24492 3936
rect 24544 3884 24550 3936
rect 25682 3884 25688 3936
rect 25740 3884 25746 3936
rect 27246 3884 27252 3936
rect 27304 3924 27310 3936
rect 27525 3927 27583 3933
rect 27525 3924 27537 3927
rect 27304 3896 27537 3924
rect 27304 3884 27310 3896
rect 27525 3893 27537 3896
rect 27571 3893 27583 3927
rect 27525 3887 27583 3893
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 27985 3927 28043 3933
rect 27985 3924 27997 3927
rect 27764 3896 27997 3924
rect 27764 3884 27770 3896
rect 27985 3893 27997 3896
rect 28031 3893 28043 3927
rect 28092 3924 28120 4032
rect 28258 3952 28264 4004
rect 28316 3992 28322 4004
rect 28368 3992 28396 4091
rect 28718 4088 28724 4100
rect 28776 4088 28782 4140
rect 28626 4020 28632 4072
rect 28684 4020 28690 4072
rect 28828 3992 28856 4168
rect 30006 4156 30012 4168
rect 30064 4156 30070 4208
rect 32968 4196 32996 4236
rect 35158 4224 35164 4236
rect 35216 4224 35222 4276
rect 35345 4267 35403 4273
rect 35345 4233 35357 4267
rect 35391 4264 35403 4267
rect 35802 4264 35808 4276
rect 35391 4236 35808 4264
rect 35391 4233 35403 4236
rect 35345 4227 35403 4233
rect 35802 4224 35808 4236
rect 35860 4224 35866 4276
rect 35986 4224 35992 4276
rect 36044 4264 36050 4276
rect 36541 4267 36599 4273
rect 36541 4264 36553 4267
rect 36044 4236 36553 4264
rect 36044 4224 36050 4236
rect 36541 4233 36553 4236
rect 36587 4233 36599 4267
rect 36541 4227 36599 4233
rect 30958 4168 32996 4196
rect 33594 4156 33600 4208
rect 33652 4156 33658 4208
rect 35434 4156 35440 4208
rect 35492 4156 35498 4208
rect 35618 4156 35624 4208
rect 35676 4196 35682 4208
rect 36633 4199 36691 4205
rect 36633 4196 36645 4199
rect 35676 4168 36645 4196
rect 35676 4156 35682 4168
rect 36633 4165 36645 4168
rect 36679 4165 36691 4199
rect 36633 4159 36691 4165
rect 32030 4088 32036 4140
rect 32088 4128 32094 4140
rect 32309 4131 32367 4137
rect 32309 4128 32321 4131
rect 32088 4100 32321 4128
rect 32088 4088 32094 4100
rect 32309 4097 32321 4100
rect 32355 4097 32367 4131
rect 32309 4091 32367 4097
rect 37274 4088 37280 4140
rect 37332 4128 37338 4140
rect 37461 4131 37519 4137
rect 37461 4128 37473 4131
rect 37332 4100 37473 4128
rect 37332 4088 37338 4100
rect 37461 4097 37473 4100
rect 37507 4128 37519 4131
rect 38102 4128 38108 4140
rect 37507 4100 38108 4128
rect 37507 4097 37519 4100
rect 37461 4091 37519 4097
rect 38102 4088 38108 4100
rect 38160 4088 38166 4140
rect 29454 4020 29460 4072
rect 29512 4020 29518 4072
rect 29733 4063 29791 4069
rect 29733 4029 29745 4063
rect 29779 4060 29791 4063
rect 30374 4060 30380 4072
rect 29779 4032 30380 4060
rect 29779 4029 29791 4032
rect 29733 4023 29791 4029
rect 30374 4020 30380 4032
rect 30432 4020 30438 4072
rect 32585 4063 32643 4069
rect 32585 4029 32597 4063
rect 32631 4060 32643 4063
rect 32674 4060 32680 4072
rect 32631 4032 32680 4060
rect 32631 4029 32643 4032
rect 32585 4023 32643 4029
rect 32674 4020 32680 4032
rect 32732 4020 32738 4072
rect 32950 4020 32956 4072
rect 33008 4060 33014 4072
rect 33008 4032 34560 4060
rect 33008 4020 33014 4032
rect 32122 3992 32128 4004
rect 28316 3964 28856 3992
rect 30760 3964 32128 3992
rect 28316 3952 28322 3964
rect 30760 3924 30788 3964
rect 32122 3952 32128 3964
rect 32180 3952 32186 4004
rect 34532 3992 34560 4032
rect 34974 4020 34980 4072
rect 35032 4060 35038 4072
rect 35529 4063 35587 4069
rect 35529 4060 35541 4063
rect 35032 4032 35541 4060
rect 35032 4020 35038 4032
rect 35529 4029 35541 4032
rect 35575 4060 35587 4063
rect 36725 4063 36783 4069
rect 36725 4060 36737 4063
rect 35575 4032 36737 4060
rect 35575 4029 35587 4032
rect 35529 4023 35587 4029
rect 36725 4029 36737 4032
rect 36771 4029 36783 4063
rect 36725 4023 36783 4029
rect 34532 3964 36216 3992
rect 28092 3896 30788 3924
rect 27985 3887 28043 3893
rect 30834 3884 30840 3936
rect 30892 3924 30898 3936
rect 31205 3927 31263 3933
rect 31205 3924 31217 3927
rect 30892 3896 31217 3924
rect 30892 3884 30898 3896
rect 31205 3893 31217 3896
rect 31251 3893 31263 3927
rect 31205 3887 31263 3893
rect 33134 3884 33140 3936
rect 33192 3924 33198 3936
rect 34057 3927 34115 3933
rect 34057 3924 34069 3927
rect 33192 3896 34069 3924
rect 33192 3884 33198 3896
rect 34057 3893 34069 3896
rect 34103 3893 34115 3927
rect 34057 3887 34115 3893
rect 34977 3927 35035 3933
rect 34977 3893 34989 3927
rect 35023 3924 35035 3927
rect 36078 3924 36084 3936
rect 35023 3896 36084 3924
rect 35023 3893 35035 3896
rect 34977 3887 35035 3893
rect 36078 3884 36084 3896
rect 36136 3884 36142 3936
rect 36188 3933 36216 3964
rect 36262 3952 36268 4004
rect 36320 3992 36326 4004
rect 37553 3995 37611 4001
rect 37553 3992 37565 3995
rect 36320 3964 37565 3992
rect 36320 3952 36326 3964
rect 37553 3961 37565 3964
rect 37599 3961 37611 3995
rect 37553 3955 37611 3961
rect 36173 3927 36231 3933
rect 36173 3893 36185 3927
rect 36219 3893 36231 3927
rect 36173 3887 36231 3893
rect 38194 3884 38200 3936
rect 38252 3884 38258 3936
rect 1104 3834 39192 3856
rect 1104 3782 5711 3834
rect 5763 3782 5775 3834
rect 5827 3782 5839 3834
rect 5891 3782 5903 3834
rect 5955 3782 5967 3834
rect 6019 3782 15233 3834
rect 15285 3782 15297 3834
rect 15349 3782 15361 3834
rect 15413 3782 15425 3834
rect 15477 3782 15489 3834
rect 15541 3782 24755 3834
rect 24807 3782 24819 3834
rect 24871 3782 24883 3834
rect 24935 3782 24947 3834
rect 24999 3782 25011 3834
rect 25063 3782 34277 3834
rect 34329 3782 34341 3834
rect 34393 3782 34405 3834
rect 34457 3782 34469 3834
rect 34521 3782 34533 3834
rect 34585 3782 39192 3834
rect 1104 3760 39192 3782
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2648 3692 2697 3720
rect 2648 3680 2654 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 3970 3680 3976 3732
rect 4028 3680 4034 3732
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 12158 3720 12164 3732
rect 8260 3692 12164 3720
rect 8260 3680 8266 3692
rect 12158 3680 12164 3692
rect 12216 3720 12222 3732
rect 13633 3723 13691 3729
rect 12216 3692 13584 3720
rect 12216 3680 12222 3692
rect 1670 3612 1676 3664
rect 1728 3652 1734 3664
rect 5537 3655 5595 3661
rect 1728 3624 5396 3652
rect 1728 3612 1734 3624
rect 1854 3544 1860 3596
rect 1912 3544 1918 3596
rect 3329 3587 3387 3593
rect 3329 3553 3341 3587
rect 3375 3584 3387 3587
rect 3510 3584 3516 3596
rect 3375 3556 3516 3584
rect 3375 3553 3387 3556
rect 3329 3547 3387 3553
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 4430 3544 4436 3596
rect 4488 3584 4494 3596
rect 4525 3587 4583 3593
rect 4525 3584 4537 3587
rect 4488 3556 4537 3584
rect 4488 3544 4494 3556
rect 4525 3553 4537 3556
rect 4571 3553 4583 3587
rect 4525 3547 4583 3553
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 1360 3488 1593 3516
rect 1360 3476 1366 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2832 3488 3065 3516
rect 2832 3476 2838 3488
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 4246 3516 4252 3528
rect 3191 3488 4252 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4614 3516 4620 3528
rect 4387 3488 4620 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 5368 3516 5396 3624
rect 5537 3621 5549 3655
rect 5583 3652 5595 3655
rect 6270 3652 6276 3664
rect 5583 3624 6276 3652
rect 5583 3621 5595 3624
rect 5537 3615 5595 3621
rect 6270 3612 6276 3624
rect 6328 3612 6334 3664
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 6641 3655 6699 3661
rect 6641 3652 6653 3655
rect 6604 3624 6653 3652
rect 6604 3612 6610 3624
rect 6641 3621 6653 3624
rect 6687 3621 6699 3655
rect 13556 3652 13584 3692
rect 13633 3689 13645 3723
rect 13679 3720 13691 3723
rect 13679 3692 16252 3720
rect 13679 3689 13691 3692
rect 13633 3683 13691 3689
rect 14642 3652 14648 3664
rect 13556 3624 14648 3652
rect 6641 3615 6699 3621
rect 14642 3612 14648 3624
rect 14700 3612 14706 3664
rect 16224 3652 16252 3692
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16356 3692 16681 3720
rect 16356 3680 16362 3692
rect 16669 3689 16681 3692
rect 16715 3720 16727 3723
rect 18506 3720 18512 3732
rect 16715 3692 18512 3720
rect 16715 3689 16727 3692
rect 16669 3683 16727 3689
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 18598 3680 18604 3732
rect 18656 3720 18662 3732
rect 18877 3723 18935 3729
rect 18877 3720 18889 3723
rect 18656 3692 18889 3720
rect 18656 3680 18662 3692
rect 18877 3689 18889 3692
rect 18923 3689 18935 3723
rect 19886 3720 19892 3732
rect 18877 3683 18935 3689
rect 18984 3692 19892 3720
rect 16224 3624 16712 3652
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 5994 3584 6000 3596
rect 5684 3556 6000 3584
rect 5684 3544 5690 3556
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 7098 3584 7104 3596
rect 6788 3556 7104 3584
rect 6788 3544 6794 3556
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 7282 3544 7288 3596
rect 7340 3544 7346 3596
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 8754 3584 8760 3596
rect 8527 3556 8760 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 10042 3544 10048 3596
rect 10100 3544 10106 3596
rect 10134 3544 10140 3596
rect 10192 3584 10198 3596
rect 12342 3584 12348 3596
rect 10192 3556 12348 3584
rect 10192 3544 10198 3556
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 14918 3544 14924 3596
rect 14976 3544 14982 3596
rect 15197 3587 15255 3593
rect 15197 3553 15209 3587
rect 15243 3584 15255 3587
rect 16574 3584 16580 3596
rect 15243 3556 16580 3584
rect 15243 3553 15255 3556
rect 15197 3547 15255 3553
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 5368 3488 7941 3516
rect 7929 3485 7941 3488
rect 7975 3516 7987 3519
rect 8386 3516 8392 3528
rect 7975 3488 8392 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 9861 3519 9919 3525
rect 9861 3485 9873 3519
rect 9907 3516 9919 3519
rect 11054 3516 11060 3528
rect 9907 3488 11060 3516
rect 9907 3485 9919 3488
rect 9861 3479 9919 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11330 3476 11336 3528
rect 11388 3476 11394 3528
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13044 3488 13553 3516
rect 13044 3476 13050 3488
rect 13541 3485 13553 3488
rect 13587 3516 13599 3519
rect 13814 3516 13820 3528
rect 13587 3488 13820 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 14090 3476 14096 3528
rect 14148 3516 14154 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14148 3488 14289 3516
rect 14148 3476 14154 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 16684 3516 16712 3624
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 17126 3584 17132 3596
rect 16908 3556 17132 3584
rect 16908 3544 16914 3556
rect 17126 3544 17132 3556
rect 17184 3544 17190 3596
rect 17770 3544 17776 3596
rect 17828 3584 17834 3596
rect 18984 3584 19012 3692
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 22373 3723 22431 3729
rect 20916 3692 22232 3720
rect 17828 3556 19012 3584
rect 17828 3544 17834 3556
rect 19426 3544 19432 3596
rect 19484 3544 19490 3596
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3584 19763 3587
rect 20916 3584 20944 3692
rect 21177 3655 21235 3661
rect 21177 3621 21189 3655
rect 21223 3652 21235 3655
rect 22204 3652 22232 3692
rect 22373 3689 22385 3723
rect 22419 3720 22431 3723
rect 22554 3720 22560 3732
rect 22419 3692 22560 3720
rect 22419 3689 22431 3692
rect 22373 3683 22431 3689
rect 22554 3680 22560 3692
rect 22612 3680 22618 3732
rect 25682 3720 25688 3732
rect 22664 3692 25688 3720
rect 22664 3652 22692 3692
rect 25682 3680 25688 3692
rect 25740 3680 25746 3732
rect 27249 3723 27307 3729
rect 27249 3689 27261 3723
rect 27295 3720 27307 3723
rect 27338 3720 27344 3732
rect 27295 3692 27344 3720
rect 27295 3689 27307 3692
rect 27249 3683 27307 3689
rect 27338 3680 27344 3692
rect 27396 3680 27402 3732
rect 27430 3680 27436 3732
rect 27488 3680 27494 3732
rect 28350 3680 28356 3732
rect 28408 3720 28414 3732
rect 28902 3720 28908 3732
rect 28408 3692 28908 3720
rect 28408 3680 28414 3692
rect 28902 3680 28908 3692
rect 28960 3680 28966 3732
rect 28994 3680 29000 3732
rect 29052 3720 29058 3732
rect 29917 3723 29975 3729
rect 29917 3720 29929 3723
rect 29052 3692 29929 3720
rect 29052 3680 29058 3692
rect 29917 3689 29929 3692
rect 29963 3689 29975 3723
rect 29917 3683 29975 3689
rect 30824 3723 30882 3729
rect 30824 3689 30836 3723
rect 30870 3720 30882 3723
rect 32953 3723 33011 3729
rect 32953 3720 32965 3723
rect 30870 3692 32965 3720
rect 30870 3689 30882 3692
rect 30824 3683 30882 3689
rect 32953 3689 32965 3692
rect 32999 3689 33011 3723
rect 32953 3683 33011 3689
rect 33042 3680 33048 3732
rect 33100 3720 33106 3732
rect 37274 3720 37280 3732
rect 33100 3692 37280 3720
rect 33100 3680 33106 3692
rect 37274 3680 37280 3692
rect 37332 3680 37338 3732
rect 27985 3655 28043 3661
rect 27985 3652 27997 3655
rect 21223 3624 22094 3652
rect 22204 3624 22692 3652
rect 26528 3624 27997 3652
rect 21223 3621 21235 3624
rect 21177 3615 21235 3621
rect 19751 3556 20944 3584
rect 22066 3584 22094 3624
rect 22646 3584 22652 3596
rect 22066 3556 22652 3584
rect 19751 3553 19763 3556
rect 19705 3547 19763 3553
rect 22646 3544 22652 3556
rect 22704 3544 22710 3596
rect 22922 3544 22928 3596
rect 22980 3544 22986 3596
rect 23198 3544 23204 3596
rect 23256 3584 23262 3596
rect 23845 3587 23903 3593
rect 23256 3556 23612 3584
rect 23256 3544 23262 3556
rect 16684 3488 17080 3516
rect 14277 3479 14335 3485
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 6089 3451 6147 3457
rect 6089 3448 6101 3451
rect 2924 3420 6101 3448
rect 2924 3408 2930 3420
rect 6089 3417 6101 3420
rect 6135 3448 6147 3451
rect 9674 3448 9680 3460
rect 6135 3420 9680 3448
rect 6135 3417 6147 3420
rect 6089 3411 6147 3417
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 11606 3408 11612 3460
rect 11664 3408 11670 3460
rect 12618 3408 12624 3460
rect 12676 3408 12682 3460
rect 15470 3448 15476 3460
rect 13004 3420 15476 3448
rect 4433 3383 4491 3389
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 5166 3380 5172 3392
rect 4479 3352 5172 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 5997 3383 6055 3389
rect 5997 3349 6009 3383
rect 6043 3380 6055 3383
rect 6362 3380 6368 3392
rect 6043 3352 6368 3380
rect 6043 3349 6055 3352
rect 5997 3343 6055 3349
rect 6362 3340 6368 3352
rect 6420 3380 6426 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6420 3352 7021 3380
rect 6420 3340 6426 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7009 3343 7067 3349
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 13004 3380 13032 3420
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 16482 3448 16488 3460
rect 16422 3420 16488 3448
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 7156 3352 13032 3380
rect 7156 3340 7162 3352
rect 13078 3340 13084 3392
rect 13136 3340 13142 3392
rect 14369 3383 14427 3389
rect 14369 3349 14381 3383
rect 14415 3380 14427 3383
rect 16942 3380 16948 3392
rect 14415 3352 16948 3380
rect 14415 3349 14427 3352
rect 14369 3343 14427 3349
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 17052 3380 17080 3488
rect 20806 3476 20812 3528
rect 20864 3476 20870 3528
rect 23382 3516 23388 3528
rect 21008 3488 23388 3516
rect 17402 3408 17408 3460
rect 17460 3408 17466 3460
rect 17954 3408 17960 3460
rect 18012 3408 18018 3460
rect 19794 3448 19800 3460
rect 18708 3420 19800 3448
rect 18708 3380 18736 3420
rect 19794 3408 19800 3420
rect 19852 3408 19858 3460
rect 17052 3352 18736 3380
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 21008 3380 21036 3488
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 23584 3525 23612 3556
rect 23845 3553 23857 3587
rect 23891 3584 23903 3587
rect 24394 3584 24400 3596
rect 23891 3556 24400 3584
rect 23891 3553 23903 3556
rect 23845 3547 23903 3553
rect 24394 3544 24400 3556
rect 24452 3544 24458 3596
rect 24670 3544 24676 3596
rect 24728 3584 24734 3596
rect 24765 3587 24823 3593
rect 24765 3584 24777 3587
rect 24728 3556 24777 3584
rect 24728 3544 24734 3556
rect 24765 3553 24777 3556
rect 24811 3553 24823 3587
rect 24765 3547 24823 3553
rect 25041 3587 25099 3593
rect 25041 3553 25053 3587
rect 25087 3584 25099 3587
rect 26528 3584 26556 3624
rect 27985 3621 27997 3624
rect 28031 3621 28043 3655
rect 30101 3655 30159 3661
rect 30101 3652 30113 3655
rect 27985 3615 28043 3621
rect 28460 3624 30113 3652
rect 25087 3556 26556 3584
rect 27157 3587 27215 3593
rect 25087 3553 25099 3556
rect 25041 3547 25099 3553
rect 27157 3553 27169 3587
rect 27203 3584 27215 3587
rect 28460 3584 28488 3624
rect 30101 3621 30113 3624
rect 30147 3621 30159 3655
rect 30101 3615 30159 3621
rect 31938 3612 31944 3664
rect 31996 3652 32002 3664
rect 32309 3655 32367 3661
rect 32309 3652 32321 3655
rect 31996 3624 32321 3652
rect 31996 3612 32002 3624
rect 32309 3621 32321 3624
rect 32355 3621 32367 3655
rect 32309 3615 32367 3621
rect 27203 3556 28488 3584
rect 28629 3587 28687 3593
rect 27203 3553 27215 3556
rect 27157 3547 27215 3553
rect 28629 3553 28641 3587
rect 28675 3584 28687 3587
rect 28675 3556 28764 3584
rect 28675 3553 28687 3556
rect 28629 3547 28687 3553
rect 23569 3519 23627 3525
rect 23569 3485 23581 3519
rect 23615 3485 23627 3519
rect 24026 3516 24032 3528
rect 23569 3479 23627 3485
rect 23768 3488 24032 3516
rect 21082 3408 21088 3460
rect 21140 3448 21146 3460
rect 21729 3451 21787 3457
rect 21729 3448 21741 3451
rect 21140 3420 21741 3448
rect 21140 3408 21146 3420
rect 21729 3417 21741 3420
rect 21775 3417 21787 3451
rect 21729 3411 21787 3417
rect 22741 3451 22799 3457
rect 22741 3417 22753 3451
rect 22787 3448 22799 3451
rect 23768 3448 23796 3488
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 26142 3476 26148 3528
rect 26200 3476 26206 3528
rect 27246 3476 27252 3528
rect 27304 3476 27310 3528
rect 26602 3448 26608 3460
rect 22787 3420 23796 3448
rect 26436 3420 26608 3448
rect 22787 3417 22799 3420
rect 22741 3411 22799 3417
rect 19576 3352 21036 3380
rect 19576 3340 19582 3352
rect 21266 3340 21272 3392
rect 21324 3380 21330 3392
rect 21821 3383 21879 3389
rect 21821 3380 21833 3383
rect 21324 3352 21833 3380
rect 21324 3340 21330 3352
rect 21821 3349 21833 3352
rect 21867 3349 21879 3383
rect 21821 3343 21879 3349
rect 22833 3383 22891 3389
rect 22833 3349 22845 3383
rect 22879 3380 22891 3383
rect 26436 3380 26464 3420
rect 26602 3408 26608 3420
rect 26660 3408 26666 3460
rect 26973 3451 27031 3457
rect 26973 3417 26985 3451
rect 27019 3448 27031 3451
rect 27522 3448 27528 3460
rect 27019 3420 27528 3448
rect 27019 3417 27031 3420
rect 26973 3411 27031 3417
rect 27522 3408 27528 3420
rect 27580 3408 27586 3460
rect 28442 3448 28448 3460
rect 27816 3420 28448 3448
rect 22879 3352 26464 3380
rect 26513 3383 26571 3389
rect 22879 3349 22891 3352
rect 22833 3343 22891 3349
rect 26513 3349 26525 3383
rect 26559 3380 26571 3383
rect 27816 3380 27844 3420
rect 28442 3408 28448 3420
rect 28500 3408 28506 3460
rect 28736 3448 28764 3556
rect 29454 3544 29460 3596
rect 29512 3584 29518 3596
rect 30561 3587 30619 3593
rect 30561 3584 30573 3587
rect 29512 3556 30573 3584
rect 29512 3544 29518 3556
rect 30561 3553 30573 3556
rect 30607 3584 30619 3587
rect 32030 3584 32036 3596
rect 30607 3556 32036 3584
rect 30607 3553 30619 3556
rect 30561 3547 30619 3553
rect 32030 3544 32036 3556
rect 32088 3544 32094 3596
rect 28902 3476 28908 3528
rect 28960 3516 28966 3528
rect 29638 3516 29644 3528
rect 28960 3488 29644 3516
rect 28960 3476 28966 3488
rect 29638 3476 29644 3488
rect 29696 3476 29702 3528
rect 30098 3516 30104 3528
rect 29840 3488 30104 3516
rect 29840 3482 29868 3488
rect 29748 3457 29868 3482
rect 30098 3476 30104 3488
rect 30156 3476 30162 3528
rect 32324 3516 32352 3615
rect 36630 3612 36636 3664
rect 36688 3612 36694 3664
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 33505 3587 33563 3593
rect 33505 3584 33517 3587
rect 32456 3556 33517 3584
rect 32456 3544 32462 3556
rect 33505 3553 33517 3556
rect 33551 3553 33563 3587
rect 33505 3547 33563 3553
rect 34882 3544 34888 3596
rect 34940 3584 34946 3596
rect 35802 3584 35808 3596
rect 34940 3556 35808 3584
rect 34940 3544 34946 3556
rect 35802 3544 35808 3556
rect 35860 3544 35866 3596
rect 36998 3544 37004 3596
rect 37056 3584 37062 3596
rect 37056 3556 38516 3584
rect 37056 3544 37062 3556
rect 33321 3519 33379 3525
rect 33321 3516 33333 3519
rect 32324 3488 33333 3516
rect 33321 3485 33333 3488
rect 33367 3485 33379 3519
rect 33321 3479 33379 3485
rect 34054 3476 34060 3528
rect 34112 3516 34118 3528
rect 34149 3519 34207 3525
rect 34149 3516 34161 3519
rect 34112 3488 34161 3516
rect 34112 3476 34118 3488
rect 34149 3485 34161 3488
rect 34195 3485 34207 3519
rect 34149 3479 34207 3485
rect 37090 3476 37096 3528
rect 37148 3516 37154 3528
rect 38488 3525 38516 3556
rect 37185 3519 37243 3525
rect 37185 3516 37197 3519
rect 37148 3488 37197 3516
rect 37148 3476 37154 3488
rect 37185 3485 37197 3488
rect 37231 3485 37243 3519
rect 37185 3479 37243 3485
rect 38473 3519 38531 3525
rect 38473 3485 38485 3519
rect 38519 3485 38531 3519
rect 38473 3479 38531 3485
rect 29733 3454 29868 3457
rect 29733 3451 29791 3454
rect 28736 3420 28994 3448
rect 26559 3352 27844 3380
rect 26559 3349 26571 3352
rect 26513 3343 26571 3349
rect 28258 3340 28264 3392
rect 28316 3380 28322 3392
rect 28353 3383 28411 3389
rect 28353 3380 28365 3383
rect 28316 3352 28365 3380
rect 28316 3340 28322 3352
rect 28353 3349 28365 3352
rect 28399 3349 28411 3383
rect 28966 3380 28994 3420
rect 29733 3417 29745 3451
rect 29779 3417 29791 3451
rect 29733 3411 29791 3417
rect 29949 3451 30007 3457
rect 29949 3417 29961 3451
rect 29995 3448 30007 3451
rect 30466 3448 30472 3460
rect 29995 3420 30472 3448
rect 29995 3417 30007 3420
rect 29949 3411 30007 3417
rect 30466 3408 30472 3420
rect 30524 3408 30530 3460
rect 34790 3448 34796 3460
rect 32062 3420 34796 3448
rect 34790 3408 34796 3420
rect 34848 3408 34854 3460
rect 35158 3408 35164 3460
rect 35216 3408 35222 3460
rect 37001 3451 37059 3457
rect 37001 3448 37013 3451
rect 36386 3420 37013 3448
rect 31478 3380 31484 3392
rect 28966 3352 31484 3380
rect 28353 3343 28411 3349
rect 31478 3340 31484 3352
rect 31536 3340 31542 3392
rect 33318 3340 33324 3392
rect 33376 3380 33382 3392
rect 33413 3383 33471 3389
rect 33413 3380 33425 3383
rect 33376 3352 33425 3380
rect 33376 3340 33382 3352
rect 33413 3349 33425 3352
rect 33459 3349 33471 3383
rect 33413 3343 33471 3349
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 34241 3383 34299 3389
rect 34241 3380 34253 3383
rect 33652 3352 34253 3380
rect 33652 3340 33658 3352
rect 34241 3349 34253 3352
rect 34287 3349 34299 3383
rect 34241 3343 34299 3349
rect 35894 3340 35900 3392
rect 35952 3380 35958 3392
rect 36464 3380 36492 3420
rect 37001 3417 37013 3420
rect 37047 3417 37059 3451
rect 37001 3411 37059 3417
rect 38654 3408 38660 3460
rect 38712 3408 38718 3460
rect 35952 3352 36492 3380
rect 35952 3340 35958 3352
rect 37274 3340 37280 3392
rect 37332 3340 37338 3392
rect 1104 3290 39352 3312
rect 1104 3238 10472 3290
rect 10524 3238 10536 3290
rect 10588 3238 10600 3290
rect 10652 3238 10664 3290
rect 10716 3238 10728 3290
rect 10780 3238 19994 3290
rect 20046 3238 20058 3290
rect 20110 3238 20122 3290
rect 20174 3238 20186 3290
rect 20238 3238 20250 3290
rect 20302 3238 29516 3290
rect 29568 3238 29580 3290
rect 29632 3238 29644 3290
rect 29696 3238 29708 3290
rect 29760 3238 29772 3290
rect 29824 3238 39038 3290
rect 39090 3238 39102 3290
rect 39154 3238 39166 3290
rect 39218 3238 39230 3290
rect 39282 3238 39294 3290
rect 39346 3238 39352 3290
rect 1104 3216 39352 3238
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 5258 3176 5264 3188
rect 4663 3148 5264 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 5718 3136 5724 3188
rect 5776 3136 5782 3188
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 7377 3179 7435 3185
rect 7377 3176 7389 3179
rect 7340 3148 7389 3176
rect 7340 3136 7346 3148
rect 7377 3145 7389 3148
rect 7423 3145 7435 3179
rect 7377 3139 7435 3145
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 10321 3179 10379 3185
rect 10321 3176 10333 3179
rect 8168 3148 10333 3176
rect 8168 3136 8174 3148
rect 10321 3145 10333 3148
rect 10367 3145 10379 3179
rect 10321 3139 10379 3145
rect 11606 3136 11612 3188
rect 11664 3176 11670 3188
rect 11793 3179 11851 3185
rect 11793 3176 11805 3179
rect 11664 3148 11805 3176
rect 11664 3136 11670 3148
rect 11793 3145 11805 3148
rect 11839 3145 11851 3179
rect 11793 3139 11851 3145
rect 12158 3136 12164 3188
rect 12216 3136 12222 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 13078 3176 13084 3188
rect 12299 3148 13084 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 15381 3179 15439 3185
rect 15381 3176 15393 3179
rect 13412 3148 15393 3176
rect 13412 3136 13418 3148
rect 15381 3145 15393 3148
rect 15427 3145 15439 3179
rect 15381 3139 15439 3145
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 15528 3148 18920 3176
rect 15528 3136 15534 3148
rect 1854 3068 1860 3120
rect 1912 3068 1918 3120
rect 3418 3108 3424 3120
rect 3082 3080 3424 3108
rect 3418 3068 3424 3080
rect 3476 3068 3482 3120
rect 4154 3068 4160 3120
rect 4212 3108 4218 3120
rect 4249 3111 4307 3117
rect 4249 3108 4261 3111
rect 4212 3080 4261 3108
rect 4212 3068 4218 3080
rect 4249 3077 4261 3080
rect 4295 3077 4307 3111
rect 4249 3071 4307 3077
rect 6086 3068 6092 3120
rect 6144 3108 6150 3120
rect 6144 3080 6592 3108
rect 6144 3068 6150 3080
rect 1578 3000 1584 3052
rect 1636 3000 1642 3052
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 4065 3043 4123 3049
rect 4065 3040 4077 3043
rect 3844 3012 4077 3040
rect 3844 3000 3850 3012
rect 4065 3009 4077 3012
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4338 3000 4344 3052
rect 4396 3000 4402 3052
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 4798 3040 4804 3052
rect 4479 3012 4804 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 5718 3040 5724 3052
rect 5675 3012 5724 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 3620 2904 3648 2935
rect 3694 2932 3700 2984
rect 3752 2972 3758 2984
rect 5644 2972 5672 3003
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 6564 3049 6592 3080
rect 7650 3068 7656 3120
rect 7708 3108 7714 3120
rect 8849 3111 8907 3117
rect 8849 3108 8861 3111
rect 7708 3080 8861 3108
rect 7708 3068 7714 3080
rect 8849 3077 8861 3080
rect 8895 3077 8907 3111
rect 8849 3071 8907 3077
rect 9858 3068 9864 3120
rect 9916 3068 9922 3120
rect 10965 3111 11023 3117
rect 10965 3077 10977 3111
rect 11011 3108 11023 3111
rect 11238 3108 11244 3120
rect 11011 3080 11244 3108
rect 11011 3077 11023 3080
rect 10965 3071 11023 3077
rect 11238 3068 11244 3080
rect 11296 3068 11302 3120
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 14182 3108 14188 3120
rect 11388 3080 14188 3108
rect 11388 3068 11394 3080
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 6730 3000 6736 3052
rect 6788 3000 6794 3052
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 7616 3012 7757 3040
rect 7616 3000 7622 3012
rect 7745 3009 7757 3012
rect 7791 3040 7803 3043
rect 8202 3040 8208 3052
rect 7791 3012 8208 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 12268 3012 12940 3040
rect 3752 2944 5672 2972
rect 5905 2975 5963 2981
rect 3752 2932 3758 2944
rect 5905 2941 5917 2975
rect 5951 2972 5963 2975
rect 6086 2972 6092 2984
rect 5951 2944 6092 2972
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 7006 2972 7012 2984
rect 6196 2944 7012 2972
rect 6196 2904 6224 2944
rect 7006 2932 7012 2944
rect 7064 2972 7070 2984
rect 7837 2975 7895 2981
rect 7837 2972 7849 2975
rect 7064 2944 7849 2972
rect 7064 2932 7070 2944
rect 7837 2941 7849 2944
rect 7883 2941 7895 2975
rect 7837 2935 7895 2941
rect 7926 2932 7932 2984
rect 7984 2932 7990 2984
rect 8573 2975 8631 2981
rect 8573 2941 8585 2975
rect 8619 2941 8631 2975
rect 8573 2935 8631 2941
rect 3620 2876 6224 2904
rect 6822 2864 6828 2916
rect 6880 2904 6886 2916
rect 8588 2904 8616 2935
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 12268 2972 12296 3012
rect 8904 2944 12296 2972
rect 8904 2932 8910 2944
rect 12434 2932 12440 2984
rect 12492 2932 12498 2984
rect 12912 2972 12940 3012
rect 12986 3000 12992 3052
rect 13044 3000 13050 3052
rect 13648 3049 13676 3080
rect 14182 3068 14188 3080
rect 14240 3068 14246 3120
rect 14366 3068 14372 3120
rect 14424 3068 14430 3120
rect 18892 3117 18920 3148
rect 19886 3136 19892 3188
rect 19944 3176 19950 3188
rect 21085 3179 21143 3185
rect 21085 3176 21097 3179
rect 19944 3148 21097 3176
rect 19944 3136 19950 3148
rect 21085 3145 21097 3148
rect 21131 3145 21143 3179
rect 21085 3139 21143 3145
rect 25961 3179 26019 3185
rect 25961 3145 25973 3179
rect 26007 3176 26019 3179
rect 27062 3176 27068 3188
rect 26007 3148 27068 3176
rect 26007 3145 26019 3148
rect 25961 3139 26019 3145
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 27246 3136 27252 3188
rect 27304 3176 27310 3188
rect 27617 3179 27675 3185
rect 27617 3176 27629 3179
rect 27304 3148 27629 3176
rect 27304 3136 27310 3148
rect 27617 3145 27629 3148
rect 27663 3176 27675 3179
rect 27663 3148 31754 3176
rect 27663 3145 27675 3148
rect 27617 3139 27675 3145
rect 18877 3111 18935 3117
rect 18877 3077 18889 3111
rect 18923 3077 18935 3111
rect 18877 3071 18935 3077
rect 19610 3068 19616 3120
rect 19668 3068 19674 3120
rect 20898 3108 20904 3120
rect 20838 3080 20904 3108
rect 20898 3068 20904 3080
rect 20956 3068 20962 3120
rect 22186 3068 22192 3120
rect 22244 3108 22250 3120
rect 22281 3111 22339 3117
rect 22281 3108 22293 3111
rect 22244 3080 22293 3108
rect 22244 3068 22250 3080
rect 22281 3077 22293 3080
rect 22327 3077 22339 3111
rect 24578 3108 24584 3120
rect 22281 3071 22339 3077
rect 24228 3080 24584 3108
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 15930 3000 15936 3052
rect 15988 3000 15994 3052
rect 16850 3000 16856 3052
rect 16908 3000 16914 3052
rect 18230 3000 18236 3052
rect 18288 3000 18294 3052
rect 19334 3000 19340 3052
rect 19392 3000 19398 3052
rect 23382 3000 23388 3052
rect 23440 3000 23446 3052
rect 24228 3049 24256 3080
rect 24578 3068 24584 3080
rect 24636 3068 24642 3120
rect 26050 3108 26056 3120
rect 25714 3080 26056 3108
rect 26050 3068 26056 3080
rect 26108 3068 26114 3120
rect 26513 3111 26571 3117
rect 26513 3077 26525 3111
rect 26559 3108 26571 3111
rect 27890 3108 27896 3120
rect 26559 3080 27896 3108
rect 26559 3077 26571 3080
rect 26513 3071 26571 3077
rect 27890 3068 27896 3080
rect 27948 3068 27954 3120
rect 28994 3108 29000 3120
rect 28000 3080 29000 3108
rect 24213 3043 24271 3049
rect 24213 3009 24225 3043
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 25774 3000 25780 3052
rect 25832 3040 25838 3052
rect 26421 3043 26479 3049
rect 26421 3040 26433 3043
rect 25832 3012 26433 3040
rect 25832 3000 25838 3012
rect 26421 3009 26433 3012
rect 26467 3040 26479 3043
rect 27338 3040 27344 3052
rect 26467 3012 27344 3040
rect 26467 3009 26479 3012
rect 26421 3003 26479 3009
rect 27338 3000 27344 3012
rect 27396 3000 27402 3052
rect 27522 3000 27528 3052
rect 27580 3000 27586 3052
rect 28000 3040 28028 3080
rect 28994 3068 29000 3080
rect 29052 3068 29058 3120
rect 31726 3108 31754 3148
rect 32122 3136 32128 3188
rect 32180 3176 32186 3188
rect 33962 3176 33968 3188
rect 32180 3148 32628 3176
rect 32180 3136 32186 3148
rect 31726 3080 32352 3108
rect 27632 3012 28028 3040
rect 13909 2975 13967 2981
rect 13909 2972 13921 2975
rect 12912 2944 13921 2972
rect 13909 2941 13921 2944
rect 13955 2941 13967 2975
rect 13909 2935 13967 2941
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 16816 2944 17141 2972
rect 16816 2932 16822 2944
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 22002 2932 22008 2984
rect 22060 2932 22066 2984
rect 22738 2972 22744 2984
rect 22112 2944 22744 2972
rect 6880 2876 8616 2904
rect 6880 2864 6886 2876
rect 11146 2864 11152 2916
rect 11204 2864 11210 2916
rect 22112 2904 22140 2944
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 24118 2932 24124 2984
rect 24176 2972 24182 2984
rect 24489 2975 24547 2981
rect 24489 2972 24501 2975
rect 24176 2944 24501 2972
rect 24176 2932 24182 2944
rect 24489 2941 24501 2944
rect 24535 2941 24547 2975
rect 24489 2935 24547 2941
rect 24854 2932 24860 2984
rect 24912 2972 24918 2984
rect 27632 2972 27660 3012
rect 28074 3000 28080 3052
rect 28132 3040 28138 3052
rect 28132 3012 28672 3040
rect 28132 3000 28138 3012
rect 24912 2944 27660 2972
rect 27801 2975 27859 2981
rect 24912 2932 24918 2944
rect 27801 2941 27813 2975
rect 27847 2972 27859 2975
rect 28534 2972 28540 2984
rect 27847 2944 28540 2972
rect 27847 2941 27859 2944
rect 27801 2935 27859 2941
rect 28534 2932 28540 2944
rect 28592 2932 28598 2984
rect 28644 2981 28672 3012
rect 30006 3000 30012 3052
rect 30064 3000 30070 3052
rect 31021 3043 31079 3049
rect 31021 3040 31033 3043
rect 30116 3012 31033 3040
rect 28629 2975 28687 2981
rect 28629 2941 28641 2975
rect 28675 2941 28687 2975
rect 28629 2935 28687 2941
rect 28902 2932 28908 2984
rect 28960 2932 28966 2984
rect 20640 2876 22140 2904
rect 5261 2839 5319 2845
rect 5261 2805 5273 2839
rect 5307 2836 5319 2839
rect 6730 2836 6736 2848
rect 5307 2808 6736 2836
rect 5307 2805 5319 2808
rect 5261 2799 5319 2805
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 6914 2796 6920 2848
rect 6972 2836 6978 2848
rect 11054 2836 11060 2848
rect 6972 2808 11060 2836
rect 6972 2796 6978 2808
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 13998 2836 14004 2848
rect 13127 2808 14004 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 13998 2796 14004 2808
rect 14056 2796 14062 2848
rect 14090 2796 14096 2848
rect 14148 2836 14154 2848
rect 16025 2839 16083 2845
rect 16025 2836 16037 2839
rect 14148 2808 16037 2836
rect 14148 2796 14154 2808
rect 16025 2805 16037 2808
rect 16071 2805 16083 2839
rect 16025 2799 16083 2805
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 20640 2836 20668 2876
rect 25498 2864 25504 2916
rect 25556 2904 25562 2916
rect 27157 2907 27215 2913
rect 27157 2904 27169 2907
rect 25556 2876 27169 2904
rect 25556 2864 25562 2876
rect 27157 2873 27169 2876
rect 27203 2873 27215 2907
rect 27157 2867 27215 2873
rect 27540 2876 28764 2904
rect 19392 2808 20668 2836
rect 19392 2796 19398 2808
rect 20898 2796 20904 2848
rect 20956 2836 20962 2848
rect 23753 2839 23811 2845
rect 23753 2836 23765 2839
rect 20956 2808 23765 2836
rect 20956 2796 20962 2808
rect 23753 2805 23765 2808
rect 23799 2805 23811 2839
rect 23753 2799 23811 2805
rect 24302 2796 24308 2848
rect 24360 2836 24366 2848
rect 27540 2836 27568 2876
rect 24360 2808 27568 2836
rect 24360 2796 24366 2808
rect 27614 2796 27620 2848
rect 27672 2836 27678 2848
rect 28074 2836 28080 2848
rect 27672 2808 28080 2836
rect 27672 2796 27678 2808
rect 28074 2796 28080 2808
rect 28132 2796 28138 2848
rect 28736 2836 28764 2876
rect 30116 2848 30144 3012
rect 31021 3009 31033 3012
rect 31067 3040 31079 3043
rect 31846 3040 31852 3052
rect 31067 3012 31852 3040
rect 31067 3009 31079 3012
rect 31021 3003 31079 3009
rect 31846 3000 31852 3012
rect 31904 3000 31910 3052
rect 32324 3049 32352 3080
rect 32490 3068 32496 3120
rect 32548 3068 32554 3120
rect 32600 3117 32628 3148
rect 32692 3148 33968 3176
rect 32585 3111 32643 3117
rect 32585 3077 32597 3111
rect 32631 3077 32643 3111
rect 32585 3071 32643 3077
rect 32692 3049 32720 3148
rect 33962 3136 33968 3148
rect 34020 3136 34026 3188
rect 37458 3176 37464 3188
rect 34256 3148 37464 3176
rect 33410 3068 33416 3120
rect 33468 3068 33474 3120
rect 34256 3117 34284 3148
rect 37458 3136 37464 3148
rect 37516 3136 37522 3188
rect 34241 3111 34299 3117
rect 34241 3077 34253 3111
rect 34287 3077 34299 3111
rect 34241 3071 34299 3077
rect 34698 3068 34704 3120
rect 34756 3108 34762 3120
rect 34793 3111 34851 3117
rect 34793 3108 34805 3111
rect 34756 3080 34805 3108
rect 34756 3068 34762 3080
rect 34793 3077 34805 3080
rect 34839 3108 34851 3111
rect 34839 3080 35834 3108
rect 34839 3077 34851 3080
rect 34793 3071 34851 3077
rect 36814 3068 36820 3120
rect 36872 3108 36878 3120
rect 38473 3111 38531 3117
rect 38473 3108 38485 3111
rect 36872 3080 38485 3108
rect 36872 3068 36878 3080
rect 38473 3077 38485 3080
rect 38519 3077 38531 3111
rect 38473 3071 38531 3077
rect 32309 3043 32367 3049
rect 32309 3009 32321 3043
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 32677 3043 32735 3049
rect 32677 3009 32689 3043
rect 32723 3009 32735 3043
rect 33965 3043 34023 3049
rect 33965 3040 33977 3043
rect 32677 3003 32735 3009
rect 32876 3012 33977 3040
rect 31573 2975 31631 2981
rect 31573 2941 31585 2975
rect 31619 2972 31631 2975
rect 31864 2972 31892 3000
rect 32876 2972 32904 3012
rect 33965 3009 33977 3012
rect 34011 3009 34023 3043
rect 33965 3003 34023 3009
rect 34882 3000 34888 3052
rect 34940 3040 34946 3052
rect 35069 3043 35127 3049
rect 35069 3040 35081 3043
rect 34940 3012 35081 3040
rect 34940 3000 34946 3012
rect 35069 3009 35081 3012
rect 35115 3009 35127 3043
rect 35069 3003 35127 3009
rect 37090 3000 37096 3052
rect 37148 3040 37154 3052
rect 37461 3043 37519 3049
rect 37461 3040 37473 3043
rect 37148 3012 37473 3040
rect 37148 3000 37154 3012
rect 37461 3009 37473 3012
rect 37507 3009 37519 3043
rect 37461 3003 37519 3009
rect 31619 2944 31754 2972
rect 31864 2944 32904 2972
rect 31619 2941 31631 2944
rect 31573 2935 31631 2941
rect 30098 2836 30104 2848
rect 28736 2808 30104 2836
rect 30098 2796 30104 2808
rect 30156 2796 30162 2848
rect 30374 2796 30380 2848
rect 30432 2796 30438 2848
rect 31726 2836 31754 2944
rect 33502 2932 33508 2984
rect 33560 2932 33566 2984
rect 35345 2975 35403 2981
rect 35345 2972 35357 2975
rect 34256 2944 35357 2972
rect 32306 2864 32312 2916
rect 32364 2904 32370 2916
rect 32861 2907 32919 2913
rect 32861 2904 32873 2907
rect 32364 2876 32873 2904
rect 32364 2864 32370 2876
rect 32861 2873 32873 2876
rect 32907 2873 32919 2907
rect 33520 2904 33548 2932
rect 34256 2904 34284 2944
rect 35345 2941 35357 2944
rect 35391 2941 35403 2975
rect 35345 2935 35403 2941
rect 36814 2932 36820 2984
rect 36872 2932 36878 2984
rect 33520 2876 34284 2904
rect 38657 2907 38715 2913
rect 32861 2867 32919 2873
rect 38657 2873 38669 2907
rect 38703 2904 38715 2907
rect 39390 2904 39396 2916
rect 38703 2876 39396 2904
rect 38703 2873 38715 2876
rect 38657 2867 38715 2873
rect 39390 2864 39396 2876
rect 39448 2864 39454 2916
rect 33042 2836 33048 2848
rect 31726 2808 33048 2836
rect 33042 2796 33048 2808
rect 33100 2796 33106 2848
rect 33134 2796 33140 2848
rect 33192 2836 33198 2848
rect 33505 2839 33563 2845
rect 33505 2836 33517 2839
rect 33192 2808 33517 2836
rect 33192 2796 33198 2808
rect 33505 2805 33517 2808
rect 33551 2805 33563 2839
rect 33505 2799 33563 2805
rect 37550 2796 37556 2848
rect 37608 2796 37614 2848
rect 1104 2746 39192 2768
rect 1104 2694 5711 2746
rect 5763 2694 5775 2746
rect 5827 2694 5839 2746
rect 5891 2694 5903 2746
rect 5955 2694 5967 2746
rect 6019 2694 15233 2746
rect 15285 2694 15297 2746
rect 15349 2694 15361 2746
rect 15413 2694 15425 2746
rect 15477 2694 15489 2746
rect 15541 2694 24755 2746
rect 24807 2694 24819 2746
rect 24871 2694 24883 2746
rect 24935 2694 24947 2746
rect 24999 2694 25011 2746
rect 25063 2694 34277 2746
rect 34329 2694 34341 2746
rect 34393 2694 34405 2746
rect 34457 2694 34469 2746
rect 34521 2694 34533 2746
rect 34585 2694 39192 2746
rect 1104 2672 39192 2694
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 4985 2635 5043 2641
rect 4985 2632 4997 2635
rect 4764 2604 4997 2632
rect 4764 2592 4770 2604
rect 4985 2601 4997 2604
rect 5031 2601 5043 2635
rect 4985 2595 5043 2601
rect 5997 2635 6055 2641
rect 5997 2601 6009 2635
rect 6043 2632 6055 2635
rect 12894 2632 12900 2644
rect 6043 2604 12900 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 15838 2632 15844 2644
rect 13464 2604 15844 2632
rect 7834 2524 7840 2576
rect 7892 2564 7898 2576
rect 8297 2567 8355 2573
rect 8297 2564 8309 2567
rect 7892 2536 8309 2564
rect 7892 2524 7898 2536
rect 8297 2533 8309 2536
rect 8343 2533 8355 2567
rect 8297 2527 8355 2533
rect 9490 2524 9496 2576
rect 9548 2564 9554 2576
rect 9548 2536 11040 2564
rect 9548 2524 9554 2536
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 3602 2496 3608 2508
rect 2363 2468 3608 2496
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 5626 2496 5632 2508
rect 4448 2468 5632 2496
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 2056 2292 2084 2391
rect 2958 2388 2964 2440
rect 3016 2388 3022 2440
rect 4448 2437 4476 2468
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 6454 2496 6460 2508
rect 5736 2468 6460 2496
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2397 4491 2431
rect 4433 2391 4491 2397
rect 4798 2388 4804 2440
rect 4856 2388 4862 2440
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5736 2428 5764 2468
rect 6454 2456 6460 2468
rect 6512 2456 6518 2508
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 6822 2496 6828 2508
rect 6595 2468 6828 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 8386 2456 8392 2508
rect 8444 2496 8450 2508
rect 9861 2499 9919 2505
rect 9861 2496 9873 2499
rect 8444 2468 9873 2496
rect 8444 2456 8450 2468
rect 9861 2465 9873 2468
rect 9907 2465 9919 2499
rect 11012 2496 11040 2536
rect 11790 2524 11796 2576
rect 11848 2524 11854 2576
rect 11882 2524 11888 2576
rect 11940 2564 11946 2576
rect 12986 2564 12992 2576
rect 11940 2536 12992 2564
rect 11940 2524 11946 2536
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 12345 2499 12403 2505
rect 12345 2496 12357 2499
rect 11012 2468 12357 2496
rect 9861 2459 9919 2465
rect 12345 2465 12357 2468
rect 12391 2465 12403 2499
rect 13464 2496 13492 2604
rect 15838 2592 15844 2604
rect 15896 2592 15902 2644
rect 16025 2635 16083 2641
rect 16025 2601 16037 2635
rect 16071 2632 16083 2635
rect 17862 2632 17868 2644
rect 16071 2604 17868 2632
rect 16071 2601 16083 2604
rect 16025 2595 16083 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 18601 2635 18659 2641
rect 18601 2632 18613 2635
rect 18196 2604 18613 2632
rect 18196 2592 18202 2604
rect 18601 2601 18613 2604
rect 18647 2601 18659 2635
rect 18601 2595 18659 2601
rect 21174 2592 21180 2644
rect 21232 2592 21238 2644
rect 22544 2635 22602 2641
rect 22544 2601 22556 2635
rect 22590 2632 22602 2635
rect 24486 2632 24492 2644
rect 22590 2604 24492 2632
rect 22590 2601 22602 2604
rect 22544 2595 22602 2601
rect 24486 2592 24492 2604
rect 24544 2592 24550 2644
rect 26326 2592 26332 2644
rect 26384 2592 26390 2644
rect 26878 2592 26884 2644
rect 26936 2632 26942 2644
rect 26936 2604 28672 2632
rect 26936 2592 26942 2604
rect 23842 2524 23848 2576
rect 23900 2564 23906 2576
rect 24029 2567 24087 2573
rect 24029 2564 24041 2567
rect 23900 2536 24041 2564
rect 23900 2524 23906 2536
rect 24029 2533 24041 2536
rect 24075 2533 24087 2567
rect 28644 2564 28672 2604
rect 28718 2592 28724 2644
rect 28776 2632 28782 2644
rect 28905 2635 28963 2641
rect 28905 2632 28917 2635
rect 28776 2604 28917 2632
rect 28776 2592 28782 2604
rect 28905 2601 28917 2604
rect 28951 2601 28963 2635
rect 28905 2595 28963 2601
rect 30650 2592 30656 2644
rect 30708 2632 30714 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 30708 2604 30849 2632
rect 30708 2592 30714 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 30944 2604 33640 2632
rect 30944 2564 30972 2604
rect 28644 2536 30972 2564
rect 33612 2564 33640 2604
rect 33686 2592 33692 2644
rect 33744 2632 33750 2644
rect 34057 2635 34115 2641
rect 34057 2632 34069 2635
rect 33744 2604 34069 2632
rect 33744 2592 33750 2604
rect 34057 2601 34069 2604
rect 34103 2601 34115 2635
rect 34057 2595 34115 2601
rect 34977 2567 35035 2573
rect 34977 2564 34989 2567
rect 33612 2536 34989 2564
rect 24029 2527 24087 2533
rect 34977 2533 34989 2536
rect 35023 2533 35035 2567
rect 34977 2527 35035 2533
rect 35526 2524 35532 2576
rect 35584 2564 35590 2576
rect 35584 2536 37596 2564
rect 35584 2524 35590 2536
rect 12345 2459 12403 2465
rect 13004 2468 13492 2496
rect 5644 2400 5764 2428
rect 5813 2431 5871 2437
rect 3234 2320 3240 2372
rect 3292 2320 3298 2372
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 4617 2363 4675 2369
rect 4617 2360 4629 2363
rect 4212 2332 4629 2360
rect 4212 2320 4218 2332
rect 4617 2329 4629 2332
rect 4663 2329 4675 2363
rect 4617 2323 4675 2329
rect 4706 2320 4712 2372
rect 4764 2320 4770 2372
rect 5644 2369 5672 2400
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6178 2428 6184 2440
rect 5859 2400 6184 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 9585 2431 9643 2437
rect 8628 2400 9536 2428
rect 8628 2388 8634 2400
rect 5629 2363 5687 2369
rect 5629 2329 5641 2363
rect 5675 2329 5687 2363
rect 5629 2323 5687 2329
rect 5721 2363 5779 2369
rect 5721 2329 5733 2363
rect 5767 2360 5779 2363
rect 5767 2332 6408 2360
rect 5767 2329 5779 2332
rect 5721 2323 5779 2329
rect 5534 2292 5540 2304
rect 2056 2264 5540 2292
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 6380 2292 6408 2332
rect 6730 2320 6736 2372
rect 6788 2360 6794 2372
rect 6825 2363 6883 2369
rect 6825 2360 6837 2363
rect 6788 2332 6837 2360
rect 6788 2320 6794 2332
rect 6825 2329 6837 2332
rect 6871 2329 6883 2363
rect 8938 2360 8944 2372
rect 8050 2332 8944 2360
rect 6825 2323 6883 2329
rect 8938 2320 8944 2332
rect 8996 2320 9002 2372
rect 9508 2360 9536 2400
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 10042 2428 10048 2440
rect 9631 2400 10048 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 11882 2428 11888 2440
rect 11011 2400 11888 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 10980 2360 11008 2391
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 13004 2428 13032 2468
rect 14274 2456 14280 2508
rect 14332 2456 14338 2508
rect 16850 2456 16856 2508
rect 16908 2456 16914 2508
rect 17126 2456 17132 2508
rect 17184 2456 17190 2508
rect 17218 2456 17224 2508
rect 17276 2496 17282 2508
rect 17494 2496 17500 2508
rect 17276 2468 17500 2496
rect 17276 2456 17282 2468
rect 17494 2456 17500 2468
rect 17552 2496 17558 2508
rect 19797 2499 19855 2505
rect 19797 2496 19809 2499
rect 17552 2468 19809 2496
rect 17552 2456 17558 2468
rect 19797 2465 19809 2468
rect 19843 2465 19855 2499
rect 19797 2459 19855 2465
rect 22002 2456 22008 2508
rect 22060 2496 22066 2508
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 22060 2468 22293 2496
rect 22060 2456 22066 2468
rect 22281 2465 22293 2468
rect 22327 2496 22339 2499
rect 24578 2496 24584 2508
rect 22327 2468 24584 2496
rect 22327 2465 22339 2468
rect 22281 2459 22339 2465
rect 24578 2456 24584 2468
rect 24636 2496 24642 2508
rect 27157 2499 27215 2505
rect 27157 2496 27169 2499
rect 24636 2468 27169 2496
rect 24636 2456 24642 2468
rect 27157 2465 27169 2468
rect 27203 2496 27215 2499
rect 27522 2496 27528 2508
rect 27203 2468 27528 2496
rect 27203 2465 27215 2468
rect 27157 2459 27215 2465
rect 27522 2456 27528 2468
rect 27580 2456 27586 2508
rect 30009 2499 30067 2505
rect 30009 2465 30021 2499
rect 30055 2496 30067 2499
rect 31294 2496 31300 2508
rect 30055 2468 31300 2496
rect 30055 2465 30067 2468
rect 30009 2459 30067 2465
rect 31294 2456 31300 2468
rect 31352 2456 31358 2508
rect 31404 2468 31892 2496
rect 11992 2400 13032 2428
rect 13081 2431 13139 2437
rect 9508 2332 11008 2360
rect 8478 2292 8484 2304
rect 6380 2264 8484 2292
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 11057 2295 11115 2301
rect 11057 2261 11069 2295
rect 11103 2292 11115 2295
rect 11992 2292 12020 2400
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 12066 2320 12072 2372
rect 12124 2320 12130 2372
rect 11103 2264 12020 2292
rect 11103 2261 11115 2264
rect 11057 2255 11115 2261
rect 12158 2252 12164 2304
rect 12216 2292 12222 2304
rect 12253 2295 12311 2301
rect 12253 2292 12265 2295
rect 12216 2264 12265 2292
rect 12216 2252 12222 2264
rect 12253 2261 12265 2264
rect 12299 2261 12311 2295
rect 13096 2292 13124 2391
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 29733 2431 29791 2437
rect 29733 2397 29745 2431
rect 29779 2428 29791 2431
rect 30098 2428 30104 2440
rect 29779 2400 30104 2428
rect 29779 2397 29791 2400
rect 29733 2391 29791 2397
rect 30098 2388 30104 2400
rect 30156 2388 30162 2440
rect 30190 2388 30196 2440
rect 30248 2428 30254 2440
rect 31404 2428 31432 2468
rect 30248 2400 31432 2428
rect 31573 2431 31631 2437
rect 30248 2388 30254 2400
rect 31573 2397 31585 2431
rect 31619 2397 31631 2431
rect 31573 2391 31631 2397
rect 13170 2320 13176 2372
rect 13228 2360 13234 2372
rect 13449 2363 13507 2369
rect 13449 2360 13461 2363
rect 13228 2332 13461 2360
rect 13228 2320 13234 2332
rect 13449 2329 13461 2332
rect 13495 2329 13507 2363
rect 13449 2323 13507 2329
rect 14550 2320 14556 2372
rect 14608 2320 14614 2372
rect 15194 2320 15200 2372
rect 15252 2320 15258 2372
rect 18414 2360 18420 2372
rect 18354 2332 18420 2360
rect 18414 2320 18420 2332
rect 18472 2320 18478 2372
rect 21082 2320 21088 2372
rect 21140 2320 21146 2372
rect 24578 2360 24584 2372
rect 23782 2332 24584 2360
rect 24578 2320 24584 2332
rect 24636 2320 24642 2372
rect 24857 2363 24915 2369
rect 24857 2329 24869 2363
rect 24903 2360 24915 2363
rect 25130 2360 25136 2372
rect 24903 2332 25136 2360
rect 24903 2329 24915 2332
rect 24857 2323 24915 2329
rect 25130 2320 25136 2332
rect 25188 2320 25194 2372
rect 25314 2320 25320 2372
rect 25372 2320 25378 2372
rect 27433 2363 27491 2369
rect 27433 2329 27445 2363
rect 27479 2360 27491 2363
rect 27706 2360 27712 2372
rect 27479 2332 27712 2360
rect 27479 2329 27491 2332
rect 27433 2323 27491 2329
rect 27706 2320 27712 2332
rect 27764 2320 27770 2372
rect 29914 2360 29920 2372
rect 28658 2332 29920 2360
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 30742 2320 30748 2372
rect 30800 2320 30806 2372
rect 31588 2360 31616 2391
rect 31864 2360 31892 2468
rect 32030 2456 32036 2508
rect 32088 2496 32094 2508
rect 32309 2499 32367 2505
rect 32309 2496 32321 2499
rect 32088 2468 32321 2496
rect 32088 2456 32094 2468
rect 32309 2465 32321 2468
rect 32355 2465 32367 2499
rect 32309 2459 32367 2465
rect 32582 2456 32588 2508
rect 32640 2496 32646 2508
rect 36081 2499 36139 2505
rect 36081 2496 36093 2499
rect 32640 2468 36093 2496
rect 32640 2456 32646 2468
rect 36081 2465 36093 2468
rect 36127 2496 36139 2499
rect 36127 2468 36216 2496
rect 36127 2465 36139 2468
rect 36081 2459 36139 2465
rect 34054 2388 34060 2440
rect 34112 2428 34118 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34112 2400 34897 2428
rect 34112 2388 34118 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35345 2431 35403 2437
rect 35345 2397 35357 2431
rect 35391 2428 35403 2431
rect 35434 2428 35440 2440
rect 35391 2400 35440 2428
rect 35391 2397 35403 2400
rect 35345 2391 35403 2397
rect 35434 2388 35440 2400
rect 35492 2388 35498 2440
rect 32585 2363 32643 2369
rect 32585 2360 32597 2363
rect 31588 2332 31800 2360
rect 31864 2332 32597 2360
rect 17218 2292 17224 2304
rect 13096 2264 17224 2292
rect 12253 2255 12311 2261
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 27246 2292 27252 2304
rect 17920 2264 27252 2292
rect 17920 2252 17926 2264
rect 27246 2252 27252 2264
rect 27304 2252 27310 2304
rect 27338 2252 27344 2304
rect 27396 2292 27402 2304
rect 29270 2292 29276 2304
rect 27396 2264 29276 2292
rect 27396 2252 27402 2264
rect 29270 2252 29276 2264
rect 29328 2292 29334 2304
rect 31588 2292 31616 2332
rect 29328 2264 31616 2292
rect 29328 2252 29334 2264
rect 31662 2252 31668 2304
rect 31720 2252 31726 2304
rect 31772 2292 31800 2332
rect 32585 2329 32597 2332
rect 32631 2329 32643 2363
rect 32585 2323 32643 2329
rect 33226 2320 33232 2372
rect 33284 2320 33290 2372
rect 34146 2320 34152 2372
rect 34204 2360 34210 2372
rect 35621 2363 35679 2369
rect 35621 2360 35633 2363
rect 34204 2332 35633 2360
rect 34204 2320 34210 2332
rect 35621 2329 35633 2332
rect 35667 2360 35679 2363
rect 35710 2360 35716 2372
rect 35667 2332 35716 2360
rect 35667 2329 35679 2332
rect 35621 2323 35679 2329
rect 35710 2320 35716 2332
rect 35768 2320 35774 2372
rect 36188 2360 36216 2468
rect 37568 2437 37596 2536
rect 37553 2431 37611 2437
rect 37553 2397 37565 2431
rect 37599 2397 37611 2431
rect 37553 2391 37611 2397
rect 36541 2363 36599 2369
rect 36541 2360 36553 2363
rect 36188 2332 36553 2360
rect 36541 2329 36553 2332
rect 36587 2329 36599 2363
rect 36541 2323 36599 2329
rect 38470 2320 38476 2372
rect 38528 2320 38534 2372
rect 38654 2320 38660 2372
rect 38712 2320 38718 2372
rect 34054 2292 34060 2304
rect 31772 2264 34060 2292
rect 34054 2252 34060 2264
rect 34112 2252 34118 2304
rect 36630 2252 36636 2304
rect 36688 2252 36694 2304
rect 37642 2252 37648 2304
rect 37700 2252 37706 2304
rect 1104 2202 39352 2224
rect 1104 2150 10472 2202
rect 10524 2150 10536 2202
rect 10588 2150 10600 2202
rect 10652 2150 10664 2202
rect 10716 2150 10728 2202
rect 10780 2150 19994 2202
rect 20046 2150 20058 2202
rect 20110 2150 20122 2202
rect 20174 2150 20186 2202
rect 20238 2150 20250 2202
rect 20302 2150 29516 2202
rect 29568 2150 29580 2202
rect 29632 2150 29644 2202
rect 29696 2150 29708 2202
rect 29760 2150 29772 2202
rect 29824 2150 39038 2202
rect 39090 2150 39102 2202
rect 39154 2150 39166 2202
rect 39218 2150 39230 2202
rect 39282 2150 39294 2202
rect 39346 2150 39352 2202
rect 1104 2128 39352 2150
rect 3234 2048 3240 2100
rect 3292 2088 3298 2100
rect 13814 2088 13820 2100
rect 3292 2060 13820 2088
rect 3292 2048 3298 2060
rect 13814 2048 13820 2060
rect 13872 2048 13878 2100
rect 23198 2048 23204 2100
rect 23256 2088 23262 2100
rect 23256 2060 29868 2088
rect 23256 2048 23262 2060
rect 4706 1980 4712 2032
rect 4764 2020 4770 2032
rect 7006 2020 7012 2032
rect 4764 1992 7012 2020
rect 4764 1980 4770 1992
rect 7006 1980 7012 1992
rect 7064 1980 7070 2032
rect 12342 1980 12348 2032
rect 12400 2020 12406 2032
rect 29730 2020 29736 2032
rect 12400 1992 29736 2020
rect 12400 1980 12406 1992
rect 29730 1980 29736 1992
rect 29788 1980 29794 2032
rect 29840 2020 29868 2060
rect 29914 2048 29920 2100
rect 29972 2088 29978 2100
rect 35986 2088 35992 2100
rect 29972 2060 35992 2088
rect 29972 2048 29978 2060
rect 35986 2048 35992 2060
rect 36044 2048 36050 2100
rect 32582 2020 32588 2032
rect 29840 1992 32588 2020
rect 32582 1980 32588 1992
rect 32640 1980 32646 2032
rect 5442 1912 5448 1964
rect 5500 1952 5506 1964
rect 12158 1952 12164 1964
rect 5500 1924 12164 1952
rect 5500 1912 5506 1924
rect 12158 1912 12164 1924
rect 12216 1912 12222 1964
rect 16482 1912 16488 1964
rect 16540 1952 16546 1964
rect 37550 1952 37556 1964
rect 16540 1924 37556 1952
rect 16540 1912 16546 1924
rect 37550 1912 37556 1924
rect 37608 1912 37614 1964
rect 6086 1844 6092 1896
rect 6144 1884 6150 1896
rect 9490 1884 9496 1896
rect 6144 1856 9496 1884
rect 6144 1844 6150 1856
rect 9490 1844 9496 1856
rect 9548 1844 9554 1896
rect 13538 1844 13544 1896
rect 13596 1884 13602 1896
rect 29638 1884 29644 1896
rect 13596 1856 29644 1884
rect 13596 1844 13602 1856
rect 29638 1844 29644 1856
rect 29696 1844 29702 1896
rect 29730 1844 29736 1896
rect 29788 1884 29794 1896
rect 33502 1884 33508 1896
rect 29788 1856 33508 1884
rect 29788 1844 29794 1856
rect 33502 1844 33508 1856
rect 33560 1844 33566 1896
rect 6546 1776 6552 1828
rect 6604 1816 6610 1828
rect 16758 1816 16764 1828
rect 6604 1788 16764 1816
rect 6604 1776 6610 1788
rect 16758 1776 16764 1788
rect 16816 1776 16822 1828
rect 24578 1776 24584 1828
rect 24636 1816 24642 1828
rect 31662 1816 31668 1828
rect 24636 1788 31668 1816
rect 24636 1776 24642 1788
rect 31662 1776 31668 1788
rect 31720 1776 31726 1828
rect 12158 1708 12164 1760
rect 12216 1748 12222 1760
rect 30374 1748 30380 1760
rect 12216 1720 30380 1748
rect 12216 1708 12222 1720
rect 30374 1708 30380 1720
rect 30432 1708 30438 1760
rect 14550 1640 14556 1692
rect 14608 1680 14614 1692
rect 25498 1680 25504 1692
rect 14608 1652 25504 1680
rect 14608 1640 14614 1652
rect 25498 1640 25504 1652
rect 25556 1640 25562 1692
rect 29638 1640 29644 1692
rect 29696 1680 29702 1692
rect 33594 1680 33600 1692
rect 29696 1652 33600 1680
rect 29696 1640 29702 1652
rect 33594 1640 33600 1652
rect 33652 1640 33658 1692
rect 4062 1572 4068 1624
rect 4120 1612 4126 1624
rect 20714 1612 20720 1624
rect 4120 1584 20720 1612
rect 4120 1572 4126 1584
rect 20714 1572 20720 1584
rect 20772 1572 20778 1624
rect 8478 1504 8484 1556
rect 8536 1544 8542 1556
rect 16206 1544 16212 1556
rect 8536 1516 16212 1544
rect 8536 1504 8542 1516
rect 16206 1504 16212 1516
rect 16264 1504 16270 1556
rect 2314 1300 2320 1352
rect 2372 1340 2378 1352
rect 37366 1340 37372 1352
rect 2372 1312 37372 1340
rect 2372 1300 2378 1312
rect 37366 1300 37372 1312
rect 37424 1300 37430 1352
rect 7374 1232 7380 1284
rect 7432 1272 7438 1284
rect 38562 1272 38568 1284
rect 7432 1244 38568 1272
rect 7432 1232 7438 1244
rect 38562 1232 38568 1244
rect 38620 1232 38626 1284
rect 6270 1164 6276 1216
rect 6328 1204 6334 1216
rect 35158 1204 35164 1216
rect 6328 1176 35164 1204
rect 6328 1164 6334 1176
rect 35158 1164 35164 1176
rect 35216 1164 35222 1216
rect 11790 1096 11796 1148
rect 11848 1136 11854 1148
rect 28902 1136 28908 1148
rect 11848 1108 28908 1136
rect 11848 1096 11854 1108
rect 28902 1096 28908 1108
rect 28960 1096 28966 1148
rect 1854 960 1860 1012
rect 1912 1000 1918 1012
rect 3234 1000 3240 1012
rect 1912 972 3240 1000
rect 1912 960 1918 972
rect 3234 960 3240 972
rect 3292 960 3298 1012
rect 2958 892 2964 944
rect 3016 932 3022 944
rect 5166 932 5172 944
rect 3016 904 5172 932
rect 3016 892 3022 904
rect 5166 892 5172 904
rect 5224 892 5230 944
rect 11146 892 11152 944
rect 11204 932 11210 944
rect 15470 932 15476 944
rect 11204 904 15476 932
rect 11204 892 11210 904
rect 15470 892 15476 904
rect 15528 892 15534 944
rect 15930 892 15936 944
rect 15988 932 15994 944
rect 17402 932 17408 944
rect 15988 904 17408 932
rect 15988 892 15994 904
rect 17402 892 17408 904
rect 17460 892 17466 944
rect 21082 892 21088 944
rect 21140 932 21146 944
rect 22554 932 22560 944
rect 21140 904 22560 932
rect 21140 892 21146 904
rect 22554 892 22560 904
rect 22612 892 22618 944
rect 29638 892 29644 944
rect 29696 932 29702 944
rect 30742 932 30748 944
rect 29696 904 30748 932
rect 29696 892 29702 904
rect 30742 892 30748 904
rect 30800 892 30806 944
rect 31570 892 31576 944
rect 31628 932 31634 944
rect 33134 932 33140 944
rect 31628 904 33140 932
rect 31628 892 31634 904
rect 33134 892 33140 904
rect 33192 892 33198 944
rect 33502 892 33508 944
rect 33560 932 33566 944
rect 36630 932 36636 944
rect 33560 904 36636 932
rect 33560 892 33566 904
rect 36630 892 36636 904
rect 36688 892 36694 944
rect 36722 892 36728 944
rect 36780 932 36786 944
rect 37642 932 37648 944
rect 36780 904 37648 932
rect 36780 892 36786 904
rect 37642 892 37648 904
rect 37700 892 37706 944
rect 5534 76 5540 128
rect 5592 116 5598 128
rect 10226 116 10232 128
rect 5592 88 10232 116
rect 5592 76 5598 88
rect 10226 76 10232 88
rect 10284 76 10290 128
<< via1 >>
rect 16120 28228 16172 28280
rect 17132 28228 17184 28280
rect 2320 26800 2372 26852
rect 23756 26800 23808 26852
rect 26884 26732 26936 26784
rect 34152 26732 34204 26784
rect 5711 26630 5763 26682
rect 5775 26630 5827 26682
rect 5839 26630 5891 26682
rect 5903 26630 5955 26682
rect 5967 26630 6019 26682
rect 15233 26630 15285 26682
rect 15297 26630 15349 26682
rect 15361 26630 15413 26682
rect 15425 26630 15477 26682
rect 15489 26630 15541 26682
rect 24755 26630 24807 26682
rect 24819 26630 24871 26682
rect 24883 26630 24935 26682
rect 24947 26630 24999 26682
rect 25011 26630 25063 26682
rect 34277 26630 34329 26682
rect 34341 26630 34393 26682
rect 34405 26630 34457 26682
rect 34469 26630 34521 26682
rect 34533 26630 34585 26682
rect 664 26528 716 26580
rect 8024 26571 8076 26580
rect 8024 26537 8033 26571
rect 8033 26537 8067 26571
rect 8067 26537 8076 26571
rect 8024 26528 8076 26537
rect 26884 26528 26936 26580
rect 27344 26571 27396 26580
rect 27344 26537 27353 26571
rect 27353 26537 27387 26571
rect 27387 26537 27396 26571
rect 27344 26528 27396 26537
rect 27436 26528 27488 26580
rect 32496 26571 32548 26580
rect 32496 26537 32505 26571
rect 32505 26537 32539 26571
rect 32539 26537 32548 26571
rect 32496 26528 32548 26537
rect 33600 26528 33652 26580
rect 37648 26571 37700 26580
rect 37648 26537 37657 26571
rect 37657 26537 37691 26571
rect 37691 26537 37700 26571
rect 37648 26528 37700 26537
rect 15568 26460 15620 26512
rect 2320 26435 2372 26444
rect 2320 26401 2329 26435
rect 2329 26401 2363 26435
rect 2363 26401 2372 26435
rect 2320 26392 2372 26401
rect 13084 26392 13136 26444
rect 16120 26460 16172 26512
rect 2044 26367 2096 26376
rect 2044 26333 2053 26367
rect 2053 26333 2087 26367
rect 2087 26333 2096 26367
rect 2044 26324 2096 26333
rect 3976 26367 4028 26376
rect 3976 26333 3985 26367
rect 3985 26333 4019 26367
rect 4019 26333 4028 26367
rect 3976 26324 4028 26333
rect 6092 26324 6144 26376
rect 9128 26367 9180 26376
rect 9128 26333 9137 26367
rect 9137 26333 9171 26367
rect 9171 26333 9180 26367
rect 9128 26324 9180 26333
rect 11336 26324 11388 26376
rect 12992 26367 13044 26376
rect 12992 26333 13001 26367
rect 13001 26333 13035 26367
rect 13035 26333 13044 26367
rect 12992 26324 13044 26333
rect 14924 26367 14976 26376
rect 14924 26333 14933 26367
rect 14933 26333 14967 26367
rect 14967 26333 14976 26367
rect 14924 26324 14976 26333
rect 16672 26324 16724 26376
rect 17132 26367 17184 26376
rect 17132 26333 17141 26367
rect 17141 26333 17175 26367
rect 17175 26333 17184 26367
rect 17132 26324 17184 26333
rect 18144 26367 18196 26376
rect 18144 26333 18153 26367
rect 18153 26333 18187 26367
rect 18187 26333 18196 26367
rect 18144 26324 18196 26333
rect 20352 26503 20404 26512
rect 20352 26469 20361 26503
rect 20361 26469 20395 26503
rect 20395 26469 20404 26503
rect 20352 26460 20404 26469
rect 20628 26392 20680 26444
rect 22008 26367 22060 26376
rect 22008 26333 22017 26367
rect 22017 26333 22051 26367
rect 22051 26333 22060 26367
rect 22008 26324 22060 26333
rect 23296 26367 23348 26376
rect 23296 26333 23305 26367
rect 23305 26333 23339 26367
rect 23339 26333 23348 26367
rect 23296 26324 23348 26333
rect 3056 26299 3108 26308
rect 3056 26265 3065 26299
rect 3065 26265 3099 26299
rect 3099 26265 3108 26299
rect 3056 26256 3108 26265
rect 7932 26299 7984 26308
rect 7932 26265 7941 26299
rect 7941 26265 7975 26299
rect 7975 26265 7984 26299
rect 7932 26256 7984 26265
rect 9404 26299 9456 26308
rect 9404 26265 9413 26299
rect 9413 26265 9447 26299
rect 9447 26265 9456 26299
rect 9404 26256 9456 26265
rect 16948 26299 17000 26308
rect 16948 26265 16957 26299
rect 16957 26265 16991 26299
rect 16991 26265 17000 26299
rect 16948 26256 17000 26265
rect 18512 26256 18564 26308
rect 25136 26324 25188 26376
rect 23572 26299 23624 26308
rect 23572 26265 23581 26299
rect 23581 26265 23615 26299
rect 23615 26265 23624 26299
rect 23572 26256 23624 26265
rect 34704 26460 34756 26512
rect 35532 26460 35584 26512
rect 27896 26392 27948 26444
rect 11888 26231 11940 26240
rect 11888 26197 11897 26231
rect 11897 26197 11931 26231
rect 11931 26197 11940 26231
rect 11888 26188 11940 26197
rect 14924 26188 14976 26240
rect 28264 26256 28316 26308
rect 28632 26324 28684 26376
rect 29184 26435 29236 26444
rect 29184 26401 29193 26435
rect 29193 26401 29227 26435
rect 29227 26401 29236 26435
rect 29184 26392 29236 26401
rect 29000 26324 29052 26376
rect 30564 26324 30616 26376
rect 34612 26324 34664 26376
rect 36268 26367 36320 26376
rect 36268 26333 36277 26367
rect 36277 26333 36311 26367
rect 36311 26333 36320 26367
rect 36268 26324 36320 26333
rect 39396 26324 39448 26376
rect 31116 26299 31168 26308
rect 31116 26265 31125 26299
rect 31125 26265 31159 26299
rect 31159 26265 31168 26299
rect 31116 26256 31168 26265
rect 32404 26299 32456 26308
rect 32404 26265 32413 26299
rect 32413 26265 32447 26299
rect 32447 26265 32456 26299
rect 32404 26256 32456 26265
rect 37556 26299 37608 26308
rect 37556 26265 37565 26299
rect 37565 26265 37599 26299
rect 37599 26265 37608 26299
rect 37556 26256 37608 26265
rect 10472 26086 10524 26138
rect 10536 26086 10588 26138
rect 10600 26086 10652 26138
rect 10664 26086 10716 26138
rect 10728 26086 10780 26138
rect 19994 26086 20046 26138
rect 20058 26086 20110 26138
rect 20122 26086 20174 26138
rect 20186 26086 20238 26138
rect 20250 26086 20302 26138
rect 29516 26086 29568 26138
rect 29580 26086 29632 26138
rect 29644 26086 29696 26138
rect 29708 26086 29760 26138
rect 29772 26086 29824 26138
rect 39038 26086 39090 26138
rect 39102 26086 39154 26138
rect 39166 26086 39218 26138
rect 39230 26086 39282 26138
rect 39294 26086 39346 26138
rect 940 25984 992 26036
rect 18880 25984 18932 26036
rect 18144 25916 18196 25968
rect 30196 25916 30248 25968
rect 39488 25916 39540 25968
rect 2136 25848 2188 25900
rect 12992 25848 13044 25900
rect 18512 25848 18564 25900
rect 30288 25848 30340 25900
rect 37556 25891 37608 25900
rect 37556 25857 37565 25891
rect 37565 25857 37599 25891
rect 37599 25857 37608 25891
rect 37556 25848 37608 25857
rect 8392 25780 8444 25832
rect 9220 25780 9272 25832
rect 18236 25823 18288 25832
rect 18236 25789 18245 25823
rect 18245 25789 18279 25823
rect 18279 25789 18288 25823
rect 18236 25780 18288 25789
rect 14832 25712 14884 25764
rect 13820 25644 13872 25696
rect 16764 25644 16816 25696
rect 17040 25687 17092 25696
rect 17040 25653 17049 25687
rect 17049 25653 17083 25687
rect 17083 25653 17092 25687
rect 17040 25644 17092 25653
rect 17132 25644 17184 25696
rect 34888 25712 34940 25764
rect 32772 25644 32824 25696
rect 37648 25687 37700 25696
rect 37648 25653 37657 25687
rect 37657 25653 37691 25687
rect 37691 25653 37700 25687
rect 37648 25644 37700 25653
rect 37924 25644 37976 25696
rect 5711 25542 5763 25594
rect 5775 25542 5827 25594
rect 5839 25542 5891 25594
rect 5903 25542 5955 25594
rect 5967 25542 6019 25594
rect 15233 25542 15285 25594
rect 15297 25542 15349 25594
rect 15361 25542 15413 25594
rect 15425 25542 15477 25594
rect 15489 25542 15541 25594
rect 24755 25542 24807 25594
rect 24819 25542 24871 25594
rect 24883 25542 24935 25594
rect 24947 25542 24999 25594
rect 25011 25542 25063 25594
rect 34277 25542 34329 25594
rect 34341 25542 34393 25594
rect 34405 25542 34457 25594
rect 34469 25542 34521 25594
rect 34533 25542 34585 25594
rect 1032 25440 1084 25492
rect 8300 25440 8352 25492
rect 8392 25304 8444 25356
rect 17868 25304 17920 25356
rect 18236 25347 18288 25356
rect 18236 25313 18245 25347
rect 18245 25313 18279 25347
rect 18279 25313 18288 25347
rect 18236 25304 18288 25313
rect 7932 25236 7984 25288
rect 13912 25236 13964 25288
rect 18144 25236 18196 25288
rect 14832 25168 14884 25220
rect 18604 25168 18656 25220
rect 6184 25100 6236 25152
rect 7196 25143 7248 25152
rect 7196 25109 7205 25143
rect 7205 25109 7239 25143
rect 7239 25109 7248 25143
rect 7196 25100 7248 25109
rect 7656 25100 7708 25152
rect 13544 25100 13596 25152
rect 18144 25100 18196 25152
rect 20904 25440 20956 25492
rect 33324 25372 33376 25424
rect 36728 25440 36780 25492
rect 27804 25304 27856 25356
rect 30196 25304 30248 25356
rect 25136 25236 25188 25288
rect 31116 25168 31168 25220
rect 32588 25168 32640 25220
rect 28448 25100 28500 25152
rect 28816 25100 28868 25152
rect 36268 25236 36320 25288
rect 36452 25236 36504 25288
rect 36636 25236 36688 25288
rect 38936 25372 38988 25424
rect 10472 24998 10524 25050
rect 10536 24998 10588 25050
rect 10600 24998 10652 25050
rect 10664 24998 10716 25050
rect 10728 24998 10780 25050
rect 19994 24998 20046 25050
rect 20058 24998 20110 25050
rect 20122 24998 20174 25050
rect 20186 24998 20238 25050
rect 20250 24998 20302 25050
rect 29516 24998 29568 25050
rect 29580 24998 29632 25050
rect 29644 24998 29696 25050
rect 29708 24998 29760 25050
rect 29772 24998 29824 25050
rect 39038 24998 39090 25050
rect 39102 24998 39154 25050
rect 39166 24998 39218 25050
rect 39230 24998 39282 25050
rect 39294 24998 39346 25050
rect 18604 24896 18656 24948
rect 28172 24896 28224 24948
rect 30380 24896 30432 24948
rect 14096 24828 14148 24880
rect 17316 24828 17368 24880
rect 30932 24896 30984 24948
rect 34888 24896 34940 24948
rect 12256 24760 12308 24812
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 18144 24803 18196 24812
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 21640 24760 21692 24812
rect 36728 24871 36780 24880
rect 36728 24837 36737 24871
rect 36737 24837 36771 24871
rect 36771 24837 36780 24871
rect 36728 24828 36780 24837
rect 13084 24735 13136 24744
rect 13084 24701 13093 24735
rect 13093 24701 13127 24735
rect 13127 24701 13136 24735
rect 13084 24692 13136 24701
rect 13544 24692 13596 24744
rect 14740 24692 14792 24744
rect 17684 24692 17736 24744
rect 23756 24692 23808 24744
rect 23848 24735 23900 24744
rect 23848 24701 23857 24735
rect 23857 24701 23891 24735
rect 23891 24701 23900 24735
rect 23848 24692 23900 24701
rect 25504 24760 25556 24812
rect 28080 24760 28132 24812
rect 30288 24803 30340 24812
rect 30288 24769 30297 24803
rect 30297 24769 30331 24803
rect 30331 24769 30340 24803
rect 30288 24760 30340 24769
rect 31024 24760 31076 24812
rect 17408 24624 17460 24676
rect 24952 24667 25004 24676
rect 24952 24633 24961 24667
rect 24961 24633 24995 24667
rect 24995 24633 25004 24667
rect 24952 24624 25004 24633
rect 12716 24556 12768 24608
rect 14188 24556 14240 24608
rect 17040 24556 17092 24608
rect 30380 24624 30432 24676
rect 27620 24556 27672 24608
rect 31760 24692 31812 24744
rect 34152 24760 34204 24812
rect 34704 24735 34756 24744
rect 34704 24701 34713 24735
rect 34713 24701 34747 24735
rect 34747 24701 34756 24735
rect 34704 24692 34756 24701
rect 35256 24803 35308 24812
rect 35256 24769 35265 24803
rect 35265 24769 35299 24803
rect 35299 24769 35308 24803
rect 35256 24760 35308 24769
rect 36268 24760 36320 24812
rect 36544 24803 36596 24812
rect 36544 24769 36553 24803
rect 36553 24769 36587 24803
rect 36587 24769 36596 24803
rect 36544 24760 36596 24769
rect 36636 24803 36688 24812
rect 36636 24769 36645 24803
rect 36645 24769 36679 24803
rect 36679 24769 36688 24803
rect 36636 24760 36688 24769
rect 39396 24760 39448 24812
rect 35900 24692 35952 24744
rect 36084 24735 36136 24744
rect 36084 24701 36093 24735
rect 36093 24701 36127 24735
rect 36127 24701 36136 24735
rect 36084 24692 36136 24701
rect 36452 24692 36504 24744
rect 36912 24692 36964 24744
rect 38292 24735 38344 24744
rect 38292 24701 38301 24735
rect 38301 24701 38335 24735
rect 38335 24701 38344 24735
rect 38292 24692 38344 24701
rect 37648 24624 37700 24676
rect 35072 24556 35124 24608
rect 36084 24556 36136 24608
rect 5711 24454 5763 24506
rect 5775 24454 5827 24506
rect 5839 24454 5891 24506
rect 5903 24454 5955 24506
rect 5967 24454 6019 24506
rect 15233 24454 15285 24506
rect 15297 24454 15349 24506
rect 15361 24454 15413 24506
rect 15425 24454 15477 24506
rect 15489 24454 15541 24506
rect 24755 24454 24807 24506
rect 24819 24454 24871 24506
rect 24883 24454 24935 24506
rect 24947 24454 24999 24506
rect 25011 24454 25063 24506
rect 34277 24454 34329 24506
rect 34341 24454 34393 24506
rect 34405 24454 34457 24506
rect 34469 24454 34521 24506
rect 34533 24454 34585 24506
rect 8300 24395 8352 24404
rect 8300 24361 8309 24395
rect 8309 24361 8343 24395
rect 8343 24361 8352 24395
rect 8300 24352 8352 24361
rect 12440 24352 12492 24404
rect 16948 24352 17000 24404
rect 17868 24395 17920 24404
rect 17868 24361 17877 24395
rect 17877 24361 17911 24395
rect 17911 24361 17920 24395
rect 17868 24352 17920 24361
rect 28172 24395 28224 24404
rect 28172 24361 28181 24395
rect 28181 24361 28215 24395
rect 28215 24361 28224 24395
rect 28172 24352 28224 24361
rect 34704 24352 34756 24404
rect 36636 24352 36688 24404
rect 6184 24259 6236 24268
rect 6184 24225 6193 24259
rect 6193 24225 6227 24259
rect 6227 24225 6236 24259
rect 6184 24216 6236 24225
rect 6552 24216 6604 24268
rect 940 24148 992 24200
rect 11980 24216 12032 24268
rect 14740 24216 14792 24268
rect 15016 24284 15068 24336
rect 19064 24284 19116 24336
rect 17224 24216 17276 24268
rect 18144 24216 18196 24268
rect 18604 24216 18656 24268
rect 20536 24216 20588 24268
rect 34980 24259 35032 24268
rect 34980 24225 34989 24259
rect 34989 24225 35023 24259
rect 35023 24225 35032 24259
rect 34980 24216 35032 24225
rect 2228 24123 2280 24132
rect 2228 24089 2237 24123
rect 2237 24089 2271 24123
rect 2271 24089 2280 24123
rect 2228 24080 2280 24089
rect 8484 24148 8536 24200
rect 6092 24080 6144 24132
rect 6644 24080 6696 24132
rect 10324 24080 10376 24132
rect 14924 24148 14976 24200
rect 15200 24148 15252 24200
rect 15844 24191 15896 24200
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 16028 24191 16080 24200
rect 16028 24157 16037 24191
rect 16037 24157 16071 24191
rect 16071 24157 16080 24191
rect 16028 24148 16080 24157
rect 7656 24055 7708 24064
rect 7656 24021 7665 24055
rect 7665 24021 7699 24055
rect 7699 24021 7708 24055
rect 7656 24012 7708 24021
rect 8944 24012 8996 24064
rect 12624 24012 12676 24064
rect 13452 24012 13504 24064
rect 14280 24055 14332 24064
rect 14280 24021 14289 24055
rect 14289 24021 14323 24055
rect 14323 24021 14332 24055
rect 14280 24012 14332 24021
rect 14648 24055 14700 24064
rect 14648 24021 14657 24055
rect 14657 24021 14691 24055
rect 14691 24021 14700 24055
rect 14648 24012 14700 24021
rect 15108 24012 15160 24064
rect 15200 24012 15252 24064
rect 26976 24148 27028 24200
rect 23848 24080 23900 24132
rect 27712 24148 27764 24200
rect 28080 24191 28132 24200
rect 28080 24157 28089 24191
rect 28089 24157 28123 24191
rect 28123 24157 28132 24191
rect 28080 24148 28132 24157
rect 28540 24148 28592 24200
rect 32588 24191 32640 24200
rect 32588 24157 32597 24191
rect 32597 24157 32631 24191
rect 32631 24157 32640 24191
rect 32588 24148 32640 24157
rect 35072 24191 35124 24200
rect 35072 24157 35081 24191
rect 35081 24157 35115 24191
rect 35115 24157 35124 24191
rect 35072 24148 35124 24157
rect 35900 24216 35952 24268
rect 36452 24191 36504 24200
rect 36452 24157 36461 24191
rect 36461 24157 36495 24191
rect 36495 24157 36504 24191
rect 36452 24148 36504 24157
rect 36728 24148 36780 24200
rect 36912 24191 36964 24200
rect 36912 24157 36921 24191
rect 36921 24157 36955 24191
rect 36955 24157 36964 24191
rect 36912 24148 36964 24157
rect 27528 24123 27580 24132
rect 27528 24089 27537 24123
rect 27537 24089 27571 24123
rect 27571 24089 27580 24123
rect 27528 24080 27580 24089
rect 32956 24123 33008 24132
rect 32956 24089 32965 24123
rect 32965 24089 32999 24123
rect 32999 24089 33008 24123
rect 32956 24080 33008 24089
rect 19708 24012 19760 24064
rect 27620 24012 27672 24064
rect 32036 24012 32088 24064
rect 35440 24012 35492 24064
rect 37096 24055 37148 24064
rect 37096 24021 37105 24055
rect 37105 24021 37139 24055
rect 37139 24021 37148 24055
rect 37096 24012 37148 24021
rect 10472 23910 10524 23962
rect 10536 23910 10588 23962
rect 10600 23910 10652 23962
rect 10664 23910 10716 23962
rect 10728 23910 10780 23962
rect 19994 23910 20046 23962
rect 20058 23910 20110 23962
rect 20122 23910 20174 23962
rect 20186 23910 20238 23962
rect 20250 23910 20302 23962
rect 29516 23910 29568 23962
rect 29580 23910 29632 23962
rect 29644 23910 29696 23962
rect 29708 23910 29760 23962
rect 29772 23910 29824 23962
rect 39038 23910 39090 23962
rect 39102 23910 39154 23962
rect 39166 23910 39218 23962
rect 39230 23910 39282 23962
rect 39294 23910 39346 23962
rect 6644 23808 6696 23860
rect 7196 23808 7248 23860
rect 7748 23808 7800 23860
rect 12348 23808 12400 23860
rect 15568 23808 15620 23860
rect 2228 23536 2280 23588
rect 11060 23740 11112 23792
rect 4160 23672 4212 23724
rect 6920 23715 6972 23724
rect 6920 23681 6929 23715
rect 6929 23681 6963 23715
rect 6963 23681 6972 23715
rect 6920 23672 6972 23681
rect 7840 23672 7892 23724
rect 8116 23672 8168 23724
rect 4896 23604 4948 23656
rect 8208 23604 8260 23656
rect 15016 23740 15068 23792
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 13728 23672 13780 23724
rect 14004 23715 14056 23724
rect 14004 23681 14013 23715
rect 14013 23681 14047 23715
rect 14047 23681 14056 23715
rect 14004 23672 14056 23681
rect 30932 23808 30984 23860
rect 31300 23808 31352 23860
rect 16856 23672 16908 23724
rect 17316 23672 17368 23724
rect 17408 23715 17460 23724
rect 17408 23681 17417 23715
rect 17417 23681 17451 23715
rect 17451 23681 17460 23715
rect 17408 23672 17460 23681
rect 17684 23715 17736 23724
rect 17684 23681 17693 23715
rect 17693 23681 17727 23715
rect 17727 23681 17736 23715
rect 17684 23672 17736 23681
rect 25136 23740 25188 23792
rect 26424 23740 26476 23792
rect 38292 23740 38344 23792
rect 26240 23672 26292 23724
rect 30472 23672 30524 23724
rect 33048 23672 33100 23724
rect 34704 23672 34756 23724
rect 34980 23715 35032 23724
rect 34980 23681 34989 23715
rect 34989 23681 35023 23715
rect 35023 23681 35032 23715
rect 34980 23672 35032 23681
rect 35072 23672 35124 23724
rect 11520 23604 11572 23656
rect 11980 23604 12032 23656
rect 24492 23604 24544 23656
rect 29276 23604 29328 23656
rect 32956 23604 33008 23656
rect 13544 23536 13596 23588
rect 30380 23536 30432 23588
rect 2964 23468 3016 23520
rect 6828 23468 6880 23520
rect 12164 23468 12216 23520
rect 17868 23468 17920 23520
rect 26516 23468 26568 23520
rect 31852 23468 31904 23520
rect 35900 23536 35952 23588
rect 35624 23468 35676 23520
rect 5711 23366 5763 23418
rect 5775 23366 5827 23418
rect 5839 23366 5891 23418
rect 5903 23366 5955 23418
rect 5967 23366 6019 23418
rect 15233 23366 15285 23418
rect 15297 23366 15349 23418
rect 15361 23366 15413 23418
rect 15425 23366 15477 23418
rect 15489 23366 15541 23418
rect 24755 23366 24807 23418
rect 24819 23366 24871 23418
rect 24883 23366 24935 23418
rect 24947 23366 24999 23418
rect 25011 23366 25063 23418
rect 34277 23366 34329 23418
rect 34341 23366 34393 23418
rect 34405 23366 34457 23418
rect 34469 23366 34521 23418
rect 34533 23366 34585 23418
rect 8944 23264 8996 23316
rect 12440 23264 12492 23316
rect 26240 23264 26292 23316
rect 29920 23264 29972 23316
rect 2228 23196 2280 23248
rect 19156 23196 19208 23248
rect 3792 23128 3844 23180
rect 4068 23060 4120 23112
rect 4712 22992 4764 23044
rect 7012 23171 7064 23180
rect 7012 23137 7021 23171
rect 7021 23137 7055 23171
rect 7055 23137 7064 23171
rect 7012 23128 7064 23137
rect 8116 23128 8168 23180
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 11888 23060 11940 23112
rect 19248 23128 19300 23180
rect 27896 23128 27948 23180
rect 13728 23060 13780 23112
rect 14832 23060 14884 23112
rect 16672 23060 16724 23112
rect 25320 23060 25372 23112
rect 25504 23103 25556 23112
rect 25504 23069 25513 23103
rect 25513 23069 25547 23103
rect 25547 23069 25556 23103
rect 25504 23060 25556 23069
rect 11244 23035 11296 23044
rect 11244 23001 11253 23035
rect 11253 23001 11287 23035
rect 11287 23001 11296 23035
rect 11244 22992 11296 23001
rect 3516 22924 3568 22976
rect 6276 22924 6328 22976
rect 6736 22967 6788 22976
rect 6736 22933 6745 22967
rect 6745 22933 6779 22967
rect 6779 22933 6788 22967
rect 6736 22924 6788 22933
rect 9312 22967 9364 22976
rect 13544 22992 13596 23044
rect 18604 22992 18656 23044
rect 26884 22992 26936 23044
rect 33048 22992 33100 23044
rect 9312 22933 9337 22967
rect 9337 22933 9364 22967
rect 9312 22924 9364 22933
rect 13268 22924 13320 22976
rect 13452 22967 13504 22976
rect 13452 22933 13461 22967
rect 13461 22933 13495 22967
rect 13495 22933 13504 22967
rect 13452 22924 13504 22933
rect 14372 22967 14424 22976
rect 14372 22933 14381 22967
rect 14381 22933 14415 22967
rect 14415 22933 14424 22967
rect 14372 22924 14424 22933
rect 22652 22924 22704 22976
rect 24124 22924 24176 22976
rect 30012 22924 30064 22976
rect 32128 22924 32180 22976
rect 10472 22822 10524 22874
rect 10536 22822 10588 22874
rect 10600 22822 10652 22874
rect 10664 22822 10716 22874
rect 10728 22822 10780 22874
rect 19994 22822 20046 22874
rect 20058 22822 20110 22874
rect 20122 22822 20174 22874
rect 20186 22822 20238 22874
rect 20250 22822 20302 22874
rect 29516 22822 29568 22874
rect 29580 22822 29632 22874
rect 29644 22822 29696 22874
rect 29708 22822 29760 22874
rect 29772 22822 29824 22874
rect 39038 22822 39090 22874
rect 39102 22822 39154 22874
rect 39166 22822 39218 22874
rect 39230 22822 39282 22874
rect 39294 22822 39346 22874
rect 2228 22763 2280 22772
rect 2228 22729 2237 22763
rect 2237 22729 2271 22763
rect 2271 22729 2280 22763
rect 2228 22720 2280 22729
rect 9312 22720 9364 22772
rect 4068 22584 4120 22636
rect 7656 22652 7708 22704
rect 10324 22652 10376 22704
rect 18788 22720 18840 22772
rect 19064 22720 19116 22772
rect 14280 22652 14332 22704
rect 15568 22652 15620 22704
rect 17960 22652 18012 22704
rect 24400 22720 24452 22772
rect 32404 22720 32456 22772
rect 8208 22516 8260 22568
rect 8852 22516 8904 22568
rect 3976 22448 4028 22500
rect 7012 22448 7064 22500
rect 940 22380 992 22432
rect 3700 22423 3752 22432
rect 3700 22389 3709 22423
rect 3709 22389 3743 22423
rect 3743 22389 3752 22423
rect 3700 22380 3752 22389
rect 4804 22380 4856 22432
rect 5632 22380 5684 22432
rect 6184 22380 6236 22432
rect 11244 22584 11296 22636
rect 12532 22584 12584 22636
rect 13912 22627 13964 22636
rect 13912 22593 13921 22627
rect 13921 22593 13955 22627
rect 13955 22593 13964 22627
rect 13912 22584 13964 22593
rect 18420 22627 18472 22636
rect 18420 22593 18429 22627
rect 18429 22593 18463 22627
rect 18463 22593 18472 22627
rect 18420 22584 18472 22593
rect 11336 22516 11388 22568
rect 13084 22559 13136 22568
rect 13084 22525 13093 22559
rect 13093 22525 13127 22559
rect 13127 22525 13136 22559
rect 13084 22516 13136 22525
rect 14648 22516 14700 22568
rect 18696 22559 18748 22568
rect 18696 22525 18705 22559
rect 18705 22525 18739 22559
rect 18739 22525 18748 22559
rect 18696 22516 18748 22525
rect 19340 22448 19392 22500
rect 14556 22380 14608 22432
rect 28264 22652 28316 22704
rect 37096 22652 37148 22704
rect 24400 22627 24452 22636
rect 24400 22593 24409 22627
rect 24409 22593 24443 22627
rect 24443 22593 24452 22627
rect 24400 22584 24452 22593
rect 29000 22584 29052 22636
rect 31392 22627 31444 22636
rect 31392 22593 31401 22627
rect 31401 22593 31435 22627
rect 31435 22593 31444 22627
rect 31392 22584 31444 22593
rect 32956 22584 33008 22636
rect 22284 22448 22336 22500
rect 25228 22516 25280 22568
rect 26884 22516 26936 22568
rect 32128 22448 32180 22500
rect 33140 22516 33192 22568
rect 33968 22448 34020 22500
rect 5711 22278 5763 22330
rect 5775 22278 5827 22330
rect 5839 22278 5891 22330
rect 5903 22278 5955 22330
rect 5967 22278 6019 22330
rect 15233 22278 15285 22330
rect 15297 22278 15349 22330
rect 15361 22278 15413 22330
rect 15425 22278 15477 22330
rect 15489 22278 15541 22330
rect 24755 22278 24807 22330
rect 24819 22278 24871 22330
rect 24883 22278 24935 22330
rect 24947 22278 24999 22330
rect 25011 22278 25063 22330
rect 34277 22278 34329 22330
rect 34341 22278 34393 22330
rect 34405 22278 34457 22330
rect 34469 22278 34521 22330
rect 34533 22278 34585 22330
rect 4804 22176 4856 22228
rect 8944 22176 8996 22228
rect 25228 22176 25280 22228
rect 32588 22176 32640 22228
rect 3976 22108 4028 22160
rect 4896 22108 4948 22160
rect 3332 22083 3384 22092
rect 3332 22049 3341 22083
rect 3341 22049 3375 22083
rect 3375 22049 3384 22083
rect 3332 22040 3384 22049
rect 12440 22040 12492 22092
rect 13636 22108 13688 22160
rect 18604 22108 18656 22160
rect 30288 22108 30340 22160
rect 15568 22040 15620 22092
rect 17960 22040 18012 22092
rect 27712 22040 27764 22092
rect 31484 22040 31536 22092
rect 33140 22108 33192 22160
rect 13912 21972 13964 22024
rect 14832 22015 14884 22024
rect 14832 21981 14841 22015
rect 14841 21981 14875 22015
rect 14875 21981 14884 22015
rect 14832 21972 14884 21981
rect 18696 21972 18748 22024
rect 4252 21904 4304 21956
rect 3056 21879 3108 21888
rect 3056 21845 3065 21879
rect 3065 21845 3099 21879
rect 3099 21845 3108 21879
rect 3056 21836 3108 21845
rect 3608 21836 3660 21888
rect 3884 21836 3936 21888
rect 4160 21836 4212 21888
rect 4436 21879 4488 21888
rect 4436 21845 4445 21879
rect 4445 21845 4479 21879
rect 4479 21845 4488 21879
rect 4436 21836 4488 21845
rect 11704 21904 11756 21956
rect 12808 21836 12860 21888
rect 13728 21904 13780 21956
rect 18972 21904 19024 21956
rect 19248 21904 19300 21956
rect 26700 21972 26752 22024
rect 28540 22015 28592 22024
rect 28540 21981 28549 22015
rect 28549 21981 28583 22015
rect 28583 21981 28592 22015
rect 28540 21972 28592 21981
rect 28724 21972 28776 22024
rect 31024 21972 31076 22024
rect 31300 22015 31352 22024
rect 31300 21981 31309 22015
rect 31309 21981 31343 22015
rect 31343 21981 31352 22015
rect 31300 21972 31352 21981
rect 25044 21904 25096 21956
rect 12992 21836 13044 21888
rect 13360 21879 13412 21888
rect 13360 21845 13369 21879
rect 13369 21845 13403 21879
rect 13403 21845 13412 21879
rect 13360 21836 13412 21845
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 28632 21879 28684 21888
rect 28632 21845 28641 21879
rect 28641 21845 28675 21879
rect 28675 21845 28684 21879
rect 28632 21836 28684 21845
rect 29092 21836 29144 21888
rect 32772 21879 32824 21888
rect 32772 21845 32781 21879
rect 32781 21845 32815 21879
rect 32815 21845 32824 21879
rect 32772 21836 32824 21845
rect 32864 21879 32916 21888
rect 32864 21845 32873 21879
rect 32873 21845 32907 21879
rect 32907 21845 32916 21879
rect 32864 21836 32916 21845
rect 10472 21734 10524 21786
rect 10536 21734 10588 21786
rect 10600 21734 10652 21786
rect 10664 21734 10716 21786
rect 10728 21734 10780 21786
rect 19994 21734 20046 21786
rect 20058 21734 20110 21786
rect 20122 21734 20174 21786
rect 20186 21734 20238 21786
rect 20250 21734 20302 21786
rect 29516 21734 29568 21786
rect 29580 21734 29632 21786
rect 29644 21734 29696 21786
rect 29708 21734 29760 21786
rect 29772 21734 29824 21786
rect 39038 21734 39090 21786
rect 39102 21734 39154 21786
rect 39166 21734 39218 21786
rect 39230 21734 39282 21786
rect 39294 21734 39346 21786
rect 4068 21675 4120 21684
rect 4068 21641 4077 21675
rect 4077 21641 4111 21675
rect 4111 21641 4120 21675
rect 4068 21632 4120 21641
rect 4436 21632 4488 21684
rect 11980 21632 12032 21684
rect 15844 21632 15896 21684
rect 16764 21632 16816 21684
rect 4528 21496 4580 21548
rect 12624 21539 12676 21548
rect 12624 21505 12633 21539
rect 12633 21505 12667 21539
rect 12667 21505 12676 21539
rect 12624 21496 12676 21505
rect 12808 21539 12860 21548
rect 12808 21505 12817 21539
rect 12817 21505 12851 21539
rect 12851 21505 12860 21539
rect 12808 21496 12860 21505
rect 17224 21607 17276 21616
rect 17224 21573 17233 21607
rect 17233 21573 17267 21607
rect 17267 21573 17276 21607
rect 17224 21564 17276 21573
rect 27620 21632 27672 21684
rect 13176 21496 13228 21548
rect 25136 21564 25188 21616
rect 31760 21632 31812 21684
rect 28632 21564 28684 21616
rect 31392 21564 31444 21616
rect 13268 21428 13320 21480
rect 15016 21428 15068 21480
rect 16856 21428 16908 21480
rect 18972 21428 19024 21480
rect 23480 21428 23532 21480
rect 25044 21471 25096 21480
rect 25044 21437 25053 21471
rect 25053 21437 25087 21471
rect 25087 21437 25096 21471
rect 25044 21428 25096 21437
rect 19708 21360 19760 21412
rect 31024 21496 31076 21548
rect 36084 21496 36136 21548
rect 37556 21496 37608 21548
rect 28540 21471 28592 21480
rect 28540 21437 28549 21471
rect 28549 21437 28583 21471
rect 28583 21437 28592 21471
rect 28540 21428 28592 21437
rect 31300 21471 31352 21480
rect 31300 21437 31309 21471
rect 31309 21437 31343 21471
rect 31343 21437 31352 21471
rect 31300 21428 31352 21437
rect 31484 21471 31536 21480
rect 31484 21437 31493 21471
rect 31493 21437 31527 21471
rect 31527 21437 31536 21471
rect 31484 21428 31536 21437
rect 12624 21292 12676 21344
rect 30012 21335 30064 21344
rect 30012 21301 30021 21335
rect 30021 21301 30055 21335
rect 30055 21301 30064 21335
rect 30012 21292 30064 21301
rect 30840 21335 30892 21344
rect 30840 21301 30849 21335
rect 30849 21301 30883 21335
rect 30883 21301 30892 21335
rect 30840 21292 30892 21301
rect 5711 21190 5763 21242
rect 5775 21190 5827 21242
rect 5839 21190 5891 21242
rect 5903 21190 5955 21242
rect 5967 21190 6019 21242
rect 15233 21190 15285 21242
rect 15297 21190 15349 21242
rect 15361 21190 15413 21242
rect 15425 21190 15477 21242
rect 15489 21190 15541 21242
rect 24755 21190 24807 21242
rect 24819 21190 24871 21242
rect 24883 21190 24935 21242
rect 24947 21190 24999 21242
rect 25011 21190 25063 21242
rect 34277 21190 34329 21242
rect 34341 21190 34393 21242
rect 34405 21190 34457 21242
rect 34469 21190 34521 21242
rect 34533 21190 34585 21242
rect 12532 21088 12584 21140
rect 12808 21088 12860 21140
rect 23664 21088 23716 21140
rect 3056 21020 3108 21072
rect 13728 21020 13780 21072
rect 23572 21020 23624 21072
rect 27804 21131 27856 21140
rect 27804 21097 27813 21131
rect 27813 21097 27847 21131
rect 27847 21097 27856 21131
rect 27804 21088 27856 21097
rect 28724 21088 28776 21140
rect 29828 21088 29880 21140
rect 30196 21088 30248 21140
rect 6368 20952 6420 21004
rect 12624 20952 12676 21004
rect 13636 20952 13688 21004
rect 24584 20952 24636 21004
rect 25136 20995 25188 21004
rect 25136 20961 25145 20995
rect 25145 20961 25179 20995
rect 25179 20961 25188 20995
rect 25136 20952 25188 20961
rect 30840 21020 30892 21072
rect 28172 20952 28224 21004
rect 940 20884 992 20936
rect 4068 20884 4120 20936
rect 12532 20884 12584 20936
rect 13268 20927 13320 20936
rect 13268 20893 13277 20927
rect 13277 20893 13311 20927
rect 13311 20893 13320 20927
rect 13268 20884 13320 20893
rect 5540 20816 5592 20868
rect 10324 20816 10376 20868
rect 12900 20859 12952 20868
rect 12900 20825 12909 20859
rect 12909 20825 12943 20859
rect 12943 20825 12952 20859
rect 12900 20816 12952 20825
rect 12992 20816 13044 20868
rect 16672 20884 16724 20936
rect 27804 20884 27856 20936
rect 31392 20952 31444 21004
rect 33692 20952 33744 21004
rect 3976 20748 4028 20800
rect 9864 20748 9916 20800
rect 10968 20791 11020 20800
rect 10968 20757 10977 20791
rect 10977 20757 11011 20791
rect 11011 20757 11020 20791
rect 10968 20748 11020 20757
rect 13452 20748 13504 20800
rect 23572 20748 23624 20800
rect 25596 20748 25648 20800
rect 30104 20884 30156 20936
rect 31024 20927 31076 20936
rect 31024 20893 31033 20927
rect 31033 20893 31067 20927
rect 31067 20893 31076 20927
rect 31024 20884 31076 20893
rect 31760 20884 31812 20936
rect 28448 20816 28500 20868
rect 29000 20816 29052 20868
rect 28172 20791 28224 20800
rect 28172 20757 28181 20791
rect 28181 20757 28215 20791
rect 28215 20757 28224 20791
rect 28172 20748 28224 20757
rect 28264 20791 28316 20800
rect 28264 20757 28273 20791
rect 28273 20757 28307 20791
rect 28307 20757 28316 20791
rect 28264 20748 28316 20757
rect 28908 20748 28960 20800
rect 29368 20748 29420 20800
rect 29920 20791 29972 20800
rect 32864 20816 32916 20868
rect 35164 20859 35216 20868
rect 35164 20825 35173 20859
rect 35173 20825 35207 20859
rect 35207 20825 35216 20859
rect 35164 20816 35216 20825
rect 36176 20816 36228 20868
rect 38476 20859 38528 20868
rect 38476 20825 38485 20859
rect 38485 20825 38519 20859
rect 38519 20825 38528 20859
rect 38476 20816 38528 20825
rect 39396 20816 39448 20868
rect 29920 20757 29945 20791
rect 29945 20757 29972 20791
rect 29920 20748 29972 20757
rect 30932 20748 30984 20800
rect 10472 20646 10524 20698
rect 10536 20646 10588 20698
rect 10600 20646 10652 20698
rect 10664 20646 10716 20698
rect 10728 20646 10780 20698
rect 19994 20646 20046 20698
rect 20058 20646 20110 20698
rect 20122 20646 20174 20698
rect 20186 20646 20238 20698
rect 20250 20646 20302 20698
rect 29516 20646 29568 20698
rect 29580 20646 29632 20698
rect 29644 20646 29696 20698
rect 29708 20646 29760 20698
rect 29772 20646 29824 20698
rect 39038 20646 39090 20698
rect 39102 20646 39154 20698
rect 39166 20646 39218 20698
rect 39230 20646 39282 20698
rect 39294 20646 39346 20698
rect 11980 20544 12032 20596
rect 14924 20544 14976 20596
rect 15568 20544 15620 20596
rect 19800 20544 19852 20596
rect 25412 20544 25464 20596
rect 26884 20544 26936 20596
rect 28540 20544 28592 20596
rect 35164 20544 35216 20596
rect 36176 20587 36228 20596
rect 36176 20553 36185 20587
rect 36185 20553 36219 20587
rect 36219 20553 36228 20587
rect 36176 20544 36228 20553
rect 12532 20476 12584 20528
rect 12624 20476 12676 20528
rect 12900 20476 12952 20528
rect 6552 20408 6604 20460
rect 11336 20408 11388 20460
rect 22100 20476 22152 20528
rect 30012 20476 30064 20528
rect 33692 20476 33744 20528
rect 16948 20408 17000 20460
rect 21272 20408 21324 20460
rect 21916 20408 21968 20460
rect 2228 20383 2280 20392
rect 2228 20349 2237 20383
rect 2237 20349 2271 20383
rect 2271 20349 2280 20383
rect 2228 20340 2280 20349
rect 3884 20340 3936 20392
rect 11980 20340 12032 20392
rect 13268 20340 13320 20392
rect 17408 20340 17460 20392
rect 21732 20340 21784 20392
rect 23664 20451 23716 20460
rect 23664 20417 23673 20451
rect 23673 20417 23707 20451
rect 23707 20417 23716 20451
rect 23664 20408 23716 20417
rect 23848 20408 23900 20460
rect 32588 20408 32640 20460
rect 36084 20451 36136 20460
rect 36084 20417 36093 20451
rect 36093 20417 36127 20451
rect 36127 20417 36136 20451
rect 36084 20408 36136 20417
rect 23296 20340 23348 20392
rect 25504 20340 25556 20392
rect 27528 20340 27580 20392
rect 12808 20272 12860 20324
rect 13728 20272 13780 20324
rect 21088 20272 21140 20324
rect 4160 20204 4212 20256
rect 12992 20204 13044 20256
rect 13084 20204 13136 20256
rect 14924 20204 14976 20256
rect 18788 20204 18840 20256
rect 21180 20204 21232 20256
rect 22376 20204 22428 20256
rect 23112 20204 23164 20256
rect 23664 20204 23716 20256
rect 25136 20272 25188 20324
rect 29920 20340 29972 20392
rect 30288 20340 30340 20392
rect 32680 20340 32732 20392
rect 34796 20340 34848 20392
rect 25964 20204 26016 20256
rect 27160 20247 27212 20256
rect 27160 20213 27169 20247
rect 27169 20213 27203 20247
rect 27203 20213 27212 20247
rect 27160 20204 27212 20213
rect 5711 20102 5763 20154
rect 5775 20102 5827 20154
rect 5839 20102 5891 20154
rect 5903 20102 5955 20154
rect 5967 20102 6019 20154
rect 15233 20102 15285 20154
rect 15297 20102 15349 20154
rect 15361 20102 15413 20154
rect 15425 20102 15477 20154
rect 15489 20102 15541 20154
rect 24755 20102 24807 20154
rect 24819 20102 24871 20154
rect 24883 20102 24935 20154
rect 24947 20102 24999 20154
rect 25011 20102 25063 20154
rect 34277 20102 34329 20154
rect 34341 20102 34393 20154
rect 34405 20102 34457 20154
rect 34469 20102 34521 20154
rect 34533 20102 34585 20154
rect 6000 20043 6052 20052
rect 6000 20009 6009 20043
rect 6009 20009 6043 20043
rect 6043 20009 6052 20043
rect 6000 20000 6052 20009
rect 11336 20000 11388 20052
rect 13176 20000 13228 20052
rect 13912 20000 13964 20052
rect 14464 20043 14516 20052
rect 14464 20009 14473 20043
rect 14473 20009 14507 20043
rect 14507 20009 14516 20043
rect 14464 20000 14516 20009
rect 14832 20000 14884 20052
rect 4160 19932 4212 19984
rect 14556 19932 14608 19984
rect 5632 19864 5684 19916
rect 14464 19864 14516 19916
rect 22100 20000 22152 20052
rect 22192 20000 22244 20052
rect 26332 20000 26384 20052
rect 33048 20043 33100 20052
rect 33048 20009 33057 20043
rect 33057 20009 33091 20043
rect 33091 20009 33100 20043
rect 33048 20000 33100 20009
rect 20352 19932 20404 19984
rect 21180 19932 21232 19984
rect 2688 19839 2740 19848
rect 2688 19805 2697 19839
rect 2697 19805 2731 19839
rect 2731 19805 2740 19839
rect 2688 19796 2740 19805
rect 6184 19796 6236 19848
rect 11244 19796 11296 19848
rect 11612 19796 11664 19848
rect 12532 19796 12584 19848
rect 12900 19796 12952 19848
rect 13268 19796 13320 19848
rect 17684 19796 17736 19848
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 19294 19796 19346 19848
rect 21732 19864 21784 19916
rect 13636 19728 13688 19780
rect 17776 19728 17828 19780
rect 4252 19660 4304 19712
rect 4436 19660 4488 19712
rect 12808 19660 12860 19712
rect 14280 19660 14332 19712
rect 14924 19660 14976 19712
rect 17500 19660 17552 19712
rect 19248 19660 19300 19712
rect 19524 19660 19576 19712
rect 20720 19796 20772 19848
rect 21640 19839 21692 19848
rect 21640 19805 21649 19839
rect 21649 19805 21683 19839
rect 21683 19805 21692 19839
rect 21640 19796 21692 19805
rect 22376 19864 22428 19916
rect 22008 19839 22060 19848
rect 22008 19805 22017 19839
rect 22017 19805 22051 19839
rect 22051 19805 22060 19839
rect 22008 19796 22060 19805
rect 22836 19975 22888 19984
rect 22836 19941 22845 19975
rect 22845 19941 22879 19975
rect 22879 19941 22888 19975
rect 22836 19932 22888 19941
rect 31024 19796 31076 19848
rect 31668 19864 31720 19916
rect 19800 19728 19852 19780
rect 31852 19728 31904 19780
rect 32036 19728 32088 19780
rect 21824 19660 21876 19712
rect 22192 19703 22244 19712
rect 22192 19669 22201 19703
rect 22201 19669 22235 19703
rect 22235 19669 22244 19703
rect 22192 19660 22244 19669
rect 25596 19660 25648 19712
rect 36452 19660 36504 19712
rect 10472 19558 10524 19610
rect 10536 19558 10588 19610
rect 10600 19558 10652 19610
rect 10664 19558 10716 19610
rect 10728 19558 10780 19610
rect 19994 19558 20046 19610
rect 20058 19558 20110 19610
rect 20122 19558 20174 19610
rect 20186 19558 20238 19610
rect 20250 19558 20302 19610
rect 29516 19558 29568 19610
rect 29580 19558 29632 19610
rect 29644 19558 29696 19610
rect 29708 19558 29760 19610
rect 29772 19558 29824 19610
rect 39038 19558 39090 19610
rect 39102 19558 39154 19610
rect 39166 19558 39218 19610
rect 39230 19558 39282 19610
rect 39294 19558 39346 19610
rect 3884 19388 3936 19440
rect 2688 19320 2740 19372
rect 9588 19456 9640 19508
rect 13728 19456 13780 19508
rect 14004 19456 14056 19508
rect 12992 19388 13044 19440
rect 5632 19252 5684 19304
rect 5172 19184 5224 19236
rect 11336 19320 11388 19372
rect 12256 19320 12308 19372
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 13820 19320 13872 19372
rect 14280 19456 14332 19508
rect 14924 19431 14976 19440
rect 14924 19397 14933 19431
rect 14933 19397 14967 19431
rect 14967 19397 14976 19431
rect 14924 19388 14976 19397
rect 16672 19388 16724 19440
rect 19800 19388 19852 19440
rect 19892 19431 19944 19440
rect 19892 19397 19901 19431
rect 19901 19397 19935 19431
rect 19935 19397 19944 19431
rect 19892 19388 19944 19397
rect 21088 19456 21140 19508
rect 21732 19456 21784 19508
rect 22008 19456 22060 19508
rect 20444 19388 20496 19440
rect 14832 19320 14884 19372
rect 17224 19320 17276 19372
rect 18144 19320 18196 19372
rect 18788 19320 18840 19372
rect 18972 19320 19024 19372
rect 19432 19320 19484 19372
rect 20536 19320 20588 19372
rect 20720 19320 20772 19372
rect 22284 19320 22336 19372
rect 24584 19456 24636 19508
rect 24768 19456 24820 19508
rect 27528 19456 27580 19508
rect 28172 19456 28224 19508
rect 23940 19388 23992 19440
rect 30656 19388 30708 19440
rect 33140 19456 33192 19508
rect 36452 19499 36504 19508
rect 36452 19465 36461 19499
rect 36461 19465 36495 19499
rect 36495 19465 36504 19499
rect 36452 19456 36504 19465
rect 33232 19388 33284 19440
rect 33784 19388 33836 19440
rect 35900 19388 35952 19440
rect 24584 19363 24636 19372
rect 24584 19329 24593 19363
rect 24593 19329 24627 19363
rect 24627 19329 24636 19363
rect 24584 19320 24636 19329
rect 30748 19363 30800 19372
rect 30748 19329 30757 19363
rect 30757 19329 30791 19363
rect 30791 19329 30800 19363
rect 30748 19320 30800 19329
rect 30840 19320 30892 19372
rect 31116 19363 31168 19372
rect 31116 19329 31125 19363
rect 31125 19329 31159 19363
rect 31159 19329 31168 19363
rect 31116 19320 31168 19329
rect 34980 19320 35032 19372
rect 35624 19320 35676 19372
rect 12716 19295 12768 19304
rect 12716 19261 12725 19295
rect 12725 19261 12759 19295
rect 12759 19261 12768 19295
rect 12716 19252 12768 19261
rect 6000 19227 6052 19236
rect 6000 19193 6009 19227
rect 6009 19193 6043 19227
rect 6043 19193 6052 19227
rect 6000 19184 6052 19193
rect 14280 19184 14332 19236
rect 2228 19116 2280 19168
rect 6092 19116 6144 19168
rect 21180 19252 21232 19304
rect 21364 19295 21416 19304
rect 21364 19261 21373 19295
rect 21373 19261 21407 19295
rect 21407 19261 21416 19295
rect 21364 19252 21416 19261
rect 22652 19295 22704 19304
rect 22652 19261 22661 19295
rect 22661 19261 22695 19295
rect 22695 19261 22704 19295
rect 22652 19252 22704 19261
rect 27160 19252 27212 19304
rect 27896 19252 27948 19304
rect 28540 19252 28592 19304
rect 22100 19184 22152 19236
rect 20536 19116 20588 19168
rect 21180 19116 21232 19168
rect 24124 19159 24176 19168
rect 24124 19125 24133 19159
rect 24133 19125 24167 19159
rect 24167 19125 24176 19159
rect 24124 19116 24176 19125
rect 37464 19184 37516 19236
rect 34612 19116 34664 19168
rect 34704 19116 34756 19168
rect 5711 19014 5763 19066
rect 5775 19014 5827 19066
rect 5839 19014 5891 19066
rect 5903 19014 5955 19066
rect 5967 19014 6019 19066
rect 15233 19014 15285 19066
rect 15297 19014 15349 19066
rect 15361 19014 15413 19066
rect 15425 19014 15477 19066
rect 15489 19014 15541 19066
rect 24755 19014 24807 19066
rect 24819 19014 24871 19066
rect 24883 19014 24935 19066
rect 24947 19014 24999 19066
rect 25011 19014 25063 19066
rect 34277 19014 34329 19066
rect 34341 19014 34393 19066
rect 34405 19014 34457 19066
rect 34469 19014 34521 19066
rect 34533 19014 34585 19066
rect 20720 18912 20772 18964
rect 21732 18912 21784 18964
rect 26608 18912 26660 18964
rect 27804 18912 27856 18964
rect 25504 18844 25556 18896
rect 22284 18776 22336 18828
rect 25136 18776 25188 18828
rect 25412 18776 25464 18828
rect 26332 18819 26384 18828
rect 26332 18785 26341 18819
rect 26341 18785 26375 18819
rect 26375 18785 26384 18819
rect 26332 18776 26384 18785
rect 26424 18819 26476 18828
rect 26424 18785 26433 18819
rect 26433 18785 26467 18819
rect 26467 18785 26476 18819
rect 26424 18776 26476 18785
rect 4436 18708 4488 18760
rect 5632 18751 5684 18760
rect 5632 18717 5641 18751
rect 5641 18717 5675 18751
rect 5675 18717 5684 18751
rect 5632 18708 5684 18717
rect 6552 18708 6604 18760
rect 12256 18708 12308 18760
rect 19708 18708 19760 18760
rect 22744 18708 22796 18760
rect 27068 18887 27120 18896
rect 27068 18853 27077 18887
rect 27077 18853 27111 18887
rect 27111 18853 27120 18887
rect 27068 18844 27120 18853
rect 35440 18912 35492 18964
rect 26792 18776 26844 18828
rect 30656 18887 30708 18896
rect 30656 18853 30665 18887
rect 30665 18853 30699 18887
rect 30699 18853 30708 18887
rect 30656 18844 30708 18853
rect 30472 18776 30524 18828
rect 31024 18776 31076 18828
rect 33140 18776 33192 18828
rect 2872 18640 2924 18692
rect 17776 18683 17828 18692
rect 17776 18649 17785 18683
rect 17785 18649 17819 18683
rect 17819 18649 17828 18683
rect 17776 18640 17828 18649
rect 17868 18640 17920 18692
rect 19524 18640 19576 18692
rect 21088 18683 21140 18692
rect 21088 18649 21097 18683
rect 21097 18649 21131 18683
rect 21131 18649 21140 18683
rect 21088 18640 21140 18649
rect 24032 18640 24084 18692
rect 25412 18683 25464 18692
rect 25412 18649 25421 18683
rect 25421 18649 25455 18683
rect 25455 18649 25464 18683
rect 25412 18640 25464 18649
rect 28264 18708 28316 18760
rect 26884 18640 26936 18692
rect 27896 18640 27948 18692
rect 30840 18640 30892 18692
rect 31208 18683 31260 18692
rect 31208 18649 31217 18683
rect 31217 18649 31251 18683
rect 31251 18649 31260 18683
rect 31208 18640 31260 18649
rect 940 18572 992 18624
rect 5724 18615 5776 18624
rect 5724 18581 5733 18615
rect 5733 18581 5767 18615
rect 5767 18581 5776 18615
rect 5724 18572 5776 18581
rect 9036 18572 9088 18624
rect 21732 18572 21784 18624
rect 23020 18615 23072 18624
rect 23020 18581 23029 18615
rect 23029 18581 23063 18615
rect 23063 18581 23072 18615
rect 23020 18572 23072 18581
rect 23388 18615 23440 18624
rect 23388 18581 23397 18615
rect 23397 18581 23431 18615
rect 23431 18581 23440 18615
rect 23388 18572 23440 18581
rect 27160 18572 27212 18624
rect 27528 18615 27580 18624
rect 27528 18581 27537 18615
rect 27537 18581 27571 18615
rect 27571 18581 27580 18615
rect 27528 18572 27580 18581
rect 30748 18572 30800 18624
rect 31300 18572 31352 18624
rect 34060 18640 34112 18692
rect 35624 18776 35676 18828
rect 35716 18751 35768 18760
rect 35716 18717 35725 18751
rect 35725 18717 35759 18751
rect 35759 18717 35768 18751
rect 35716 18708 35768 18717
rect 37464 18819 37516 18828
rect 37464 18785 37473 18819
rect 37473 18785 37507 18819
rect 37507 18785 37516 18819
rect 37464 18776 37516 18785
rect 36820 18640 36872 18692
rect 10472 18470 10524 18522
rect 10536 18470 10588 18522
rect 10600 18470 10652 18522
rect 10664 18470 10716 18522
rect 10728 18470 10780 18522
rect 19994 18470 20046 18522
rect 20058 18470 20110 18522
rect 20122 18470 20174 18522
rect 20186 18470 20238 18522
rect 20250 18470 20302 18522
rect 29516 18470 29568 18522
rect 29580 18470 29632 18522
rect 29644 18470 29696 18522
rect 29708 18470 29760 18522
rect 29772 18470 29824 18522
rect 39038 18470 39090 18522
rect 39102 18470 39154 18522
rect 39166 18470 39218 18522
rect 39230 18470 39282 18522
rect 39294 18470 39346 18522
rect 5724 18368 5776 18420
rect 2964 18343 3016 18352
rect 2964 18309 2973 18343
rect 2973 18309 3007 18343
rect 3007 18309 3016 18343
rect 2964 18300 3016 18309
rect 3700 18300 3752 18352
rect 11244 18300 11296 18352
rect 12440 18232 12492 18284
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 2228 18164 2280 18216
rect 6920 18164 6972 18216
rect 14740 18164 14792 18216
rect 17960 18368 18012 18420
rect 19432 18368 19484 18420
rect 20628 18411 20680 18420
rect 20628 18377 20637 18411
rect 20637 18377 20671 18411
rect 20671 18377 20680 18411
rect 20628 18368 20680 18377
rect 22744 18368 22796 18420
rect 24032 18411 24084 18420
rect 24032 18377 24041 18411
rect 24041 18377 24075 18411
rect 24075 18377 24084 18411
rect 24032 18368 24084 18377
rect 24492 18368 24544 18420
rect 26516 18411 26568 18420
rect 26516 18377 26525 18411
rect 26525 18377 26559 18411
rect 26559 18377 26568 18411
rect 26516 18368 26568 18377
rect 30656 18368 30708 18420
rect 32588 18368 32640 18420
rect 37188 18368 37240 18420
rect 17500 18343 17552 18352
rect 17500 18309 17509 18343
rect 17509 18309 17543 18343
rect 17543 18309 17552 18343
rect 17500 18300 17552 18309
rect 19524 18300 19576 18352
rect 31576 18300 31628 18352
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 17868 18232 17920 18284
rect 18880 18232 18932 18284
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 19984 18232 20036 18241
rect 20536 18232 20588 18284
rect 21364 18275 21416 18284
rect 21364 18241 21373 18275
rect 21373 18241 21407 18275
rect 21407 18241 21416 18275
rect 21364 18232 21416 18241
rect 22652 18232 22704 18284
rect 22836 18232 22888 18284
rect 23204 18164 23256 18216
rect 23388 18232 23440 18284
rect 25320 18232 25372 18284
rect 25872 18275 25924 18284
rect 25872 18241 25881 18275
rect 25881 18241 25915 18275
rect 25915 18241 25924 18275
rect 25872 18232 25924 18241
rect 26608 18275 26660 18284
rect 26608 18241 26617 18275
rect 26617 18241 26651 18275
rect 26651 18241 26660 18275
rect 26608 18232 26660 18241
rect 27160 18275 27212 18284
rect 27160 18241 27169 18275
rect 27169 18241 27203 18275
rect 27203 18241 27212 18275
rect 27160 18232 27212 18241
rect 30840 18232 30892 18284
rect 31484 18232 31536 18284
rect 33968 18232 34020 18284
rect 36820 18232 36872 18284
rect 37188 18232 37240 18284
rect 23756 18164 23808 18216
rect 25136 18207 25188 18216
rect 25136 18173 25145 18207
rect 25145 18173 25179 18207
rect 25179 18173 25188 18207
rect 25136 18164 25188 18173
rect 26332 18207 26384 18216
rect 26332 18173 26341 18207
rect 26341 18173 26375 18207
rect 26375 18173 26384 18207
rect 26332 18164 26384 18173
rect 27712 18164 27764 18216
rect 31208 18164 31260 18216
rect 34152 18164 34204 18216
rect 35900 18164 35952 18216
rect 36452 18207 36504 18216
rect 36452 18173 36461 18207
rect 36461 18173 36495 18207
rect 36495 18173 36504 18207
rect 36452 18164 36504 18173
rect 26056 18096 26108 18148
rect 14924 18071 14976 18080
rect 14924 18037 14933 18071
rect 14933 18037 14967 18071
rect 14967 18037 14976 18071
rect 14924 18028 14976 18037
rect 17868 18071 17920 18080
rect 17868 18037 17877 18071
rect 17877 18037 17911 18071
rect 17911 18037 17920 18071
rect 17868 18028 17920 18037
rect 20444 18028 20496 18080
rect 26148 18071 26200 18080
rect 26148 18037 26157 18071
rect 26157 18037 26191 18071
rect 26191 18037 26200 18071
rect 26148 18028 26200 18037
rect 26976 18028 27028 18080
rect 31300 18028 31352 18080
rect 5711 17926 5763 17978
rect 5775 17926 5827 17978
rect 5839 17926 5891 17978
rect 5903 17926 5955 17978
rect 5967 17926 6019 17978
rect 15233 17926 15285 17978
rect 15297 17926 15349 17978
rect 15361 17926 15413 17978
rect 15425 17926 15477 17978
rect 15489 17926 15541 17978
rect 24755 17926 24807 17978
rect 24819 17926 24871 17978
rect 24883 17926 24935 17978
rect 24947 17926 24999 17978
rect 25011 17926 25063 17978
rect 34277 17926 34329 17978
rect 34341 17926 34393 17978
rect 34405 17926 34457 17978
rect 34469 17926 34521 17978
rect 34533 17926 34585 17978
rect 1768 17688 1820 17740
rect 22928 17824 22980 17876
rect 25780 17824 25832 17876
rect 26148 17867 26200 17876
rect 26148 17833 26157 17867
rect 26157 17833 26191 17867
rect 26191 17833 26200 17867
rect 26148 17824 26200 17833
rect 21088 17799 21140 17808
rect 21088 17765 21097 17799
rect 21097 17765 21131 17799
rect 21131 17765 21140 17799
rect 21088 17756 21140 17765
rect 27620 17824 27672 17876
rect 28724 17824 28776 17876
rect 29092 17824 29144 17876
rect 18052 17688 18104 17740
rect 2044 17663 2096 17672
rect 2044 17629 2053 17663
rect 2053 17629 2087 17663
rect 2087 17629 2096 17663
rect 2044 17620 2096 17629
rect 6644 17620 6696 17672
rect 14096 17620 14148 17672
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 20352 17620 20404 17672
rect 20536 17620 20588 17672
rect 22100 17620 22152 17672
rect 22284 17731 22336 17740
rect 22284 17697 22293 17731
rect 22293 17697 22327 17731
rect 22327 17697 22336 17731
rect 22284 17688 22336 17697
rect 17316 17552 17368 17604
rect 21088 17552 21140 17604
rect 2412 17484 2464 17536
rect 2780 17527 2832 17536
rect 2780 17493 2789 17527
rect 2789 17493 2823 17527
rect 2823 17493 2832 17527
rect 2780 17484 2832 17493
rect 17500 17484 17552 17536
rect 19800 17484 19852 17536
rect 19984 17484 20036 17536
rect 21732 17484 21784 17536
rect 23664 17620 23716 17672
rect 27160 17756 27212 17808
rect 28448 17756 28500 17808
rect 30564 17756 30616 17808
rect 32496 17756 32548 17808
rect 33968 17756 34020 17808
rect 25228 17731 25280 17740
rect 25228 17697 25237 17731
rect 25237 17697 25271 17731
rect 25271 17697 25280 17731
rect 25228 17688 25280 17697
rect 27344 17688 27396 17740
rect 31024 17731 31076 17740
rect 31024 17697 31033 17731
rect 31033 17697 31067 17731
rect 31067 17697 31076 17731
rect 31024 17688 31076 17697
rect 31300 17731 31352 17740
rect 31300 17697 31309 17731
rect 31309 17697 31343 17731
rect 31343 17697 31352 17731
rect 31300 17688 31352 17697
rect 31760 17688 31812 17740
rect 34612 17688 34664 17740
rect 35900 17688 35952 17740
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 27252 17620 27304 17672
rect 30196 17620 30248 17672
rect 30564 17620 30616 17672
rect 25964 17595 26016 17604
rect 25964 17561 25989 17595
rect 25989 17561 26016 17595
rect 25964 17552 26016 17561
rect 26884 17552 26936 17604
rect 30656 17552 30708 17604
rect 32772 17620 32824 17672
rect 33140 17620 33192 17672
rect 37188 17620 37240 17672
rect 27436 17527 27488 17536
rect 27436 17493 27445 17527
rect 27445 17493 27479 17527
rect 27479 17493 27488 17527
rect 27436 17484 27488 17493
rect 27528 17484 27580 17536
rect 30288 17484 30340 17536
rect 31208 17484 31260 17536
rect 32588 17484 32640 17536
rect 35164 17552 35216 17604
rect 10472 17382 10524 17434
rect 10536 17382 10588 17434
rect 10600 17382 10652 17434
rect 10664 17382 10716 17434
rect 10728 17382 10780 17434
rect 19994 17382 20046 17434
rect 20058 17382 20110 17434
rect 20122 17382 20174 17434
rect 20186 17382 20238 17434
rect 20250 17382 20302 17434
rect 29516 17382 29568 17434
rect 29580 17382 29632 17434
rect 29644 17382 29696 17434
rect 29708 17382 29760 17434
rect 29772 17382 29824 17434
rect 39038 17382 39090 17434
rect 39102 17382 39154 17434
rect 39166 17382 39218 17434
rect 39230 17382 39282 17434
rect 39294 17382 39346 17434
rect 6828 17280 6880 17332
rect 7380 17280 7432 17332
rect 7748 17212 7800 17264
rect 9496 17212 9548 17264
rect 13636 17280 13688 17332
rect 19800 17280 19852 17332
rect 17132 17255 17184 17264
rect 17132 17221 17141 17255
rect 17141 17221 17175 17255
rect 17175 17221 17184 17255
rect 17132 17212 17184 17221
rect 18144 17212 18196 17264
rect 23940 17323 23992 17332
rect 23940 17289 23949 17323
rect 23949 17289 23983 17323
rect 23983 17289 23992 17323
rect 23940 17280 23992 17289
rect 24124 17280 24176 17332
rect 1584 17187 1636 17196
rect 1584 17153 1593 17187
rect 1593 17153 1627 17187
rect 1627 17153 1636 17187
rect 1584 17144 1636 17153
rect 3976 17144 4028 17196
rect 5172 17187 5224 17196
rect 5172 17153 5181 17187
rect 5181 17153 5215 17187
rect 5215 17153 5224 17187
rect 5172 17144 5224 17153
rect 8024 17187 8076 17196
rect 8024 17153 8033 17187
rect 8033 17153 8067 17187
rect 8067 17153 8076 17187
rect 8024 17144 8076 17153
rect 2228 17076 2280 17128
rect 4344 17076 4396 17128
rect 5080 17008 5132 17060
rect 5540 17076 5592 17128
rect 10876 17076 10928 17128
rect 11888 17076 11940 17128
rect 13176 17144 13228 17196
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 15660 17144 15712 17196
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 1860 16940 1912 16992
rect 4436 16940 4488 16992
rect 4804 16983 4856 16992
rect 4804 16949 4813 16983
rect 4813 16949 4847 16983
rect 4847 16949 4856 16983
rect 4804 16940 4856 16949
rect 5356 16940 5408 16992
rect 6828 16940 6880 16992
rect 16488 17076 16540 17128
rect 18788 17076 18840 17128
rect 22836 17144 22888 17196
rect 20812 17076 20864 17128
rect 23388 17212 23440 17264
rect 24584 17212 24636 17264
rect 23848 17187 23900 17196
rect 23848 17153 23857 17187
rect 23857 17153 23891 17187
rect 23891 17153 23900 17187
rect 23848 17144 23900 17153
rect 24492 17187 24544 17196
rect 24492 17153 24501 17187
rect 24501 17153 24535 17187
rect 24535 17153 24544 17187
rect 24492 17144 24544 17153
rect 26332 17280 26384 17332
rect 32772 17280 32824 17332
rect 32956 17323 33008 17332
rect 32956 17289 32965 17323
rect 32965 17289 32999 17323
rect 32999 17289 33008 17323
rect 32956 17280 33008 17289
rect 26056 17187 26108 17196
rect 26056 17153 26065 17187
rect 26065 17153 26099 17187
rect 26099 17153 26108 17187
rect 26056 17144 26108 17153
rect 26700 17212 26752 17264
rect 27436 17212 27488 17264
rect 28356 17144 28408 17196
rect 29000 17144 29052 17196
rect 30104 17144 30156 17196
rect 30380 17144 30432 17196
rect 30564 17144 30616 17196
rect 30840 17187 30892 17196
rect 30840 17153 30849 17187
rect 30849 17153 30883 17187
rect 30883 17153 30892 17187
rect 30840 17144 30892 17153
rect 31024 17212 31076 17264
rect 32588 17255 32640 17264
rect 32588 17221 32597 17255
rect 32597 17221 32631 17255
rect 32631 17221 32640 17255
rect 32588 17212 32640 17221
rect 38568 17280 38620 17332
rect 33968 17212 34020 17264
rect 34336 17212 34388 17264
rect 35716 17212 35768 17264
rect 29184 17076 29236 17128
rect 29736 17076 29788 17128
rect 29920 17076 29972 17128
rect 31576 17076 31628 17128
rect 31668 17076 31720 17128
rect 21640 17008 21692 17060
rect 29368 17008 29420 17060
rect 20996 16940 21048 16992
rect 21548 16940 21600 16992
rect 27160 16940 27212 16992
rect 27620 16940 27672 16992
rect 27988 16940 28040 16992
rect 30104 16940 30156 16992
rect 30380 17008 30432 17060
rect 32680 17076 32732 17128
rect 34152 17187 34204 17196
rect 34152 17153 34161 17187
rect 34161 17153 34195 17187
rect 34195 17153 34204 17187
rect 34152 17144 34204 17153
rect 34336 17119 34388 17128
rect 34336 17085 34345 17119
rect 34345 17085 34379 17119
rect 34379 17085 34388 17119
rect 34336 17076 34388 17085
rect 34888 17144 34940 17196
rect 37372 17144 37424 17196
rect 35256 17076 35308 17128
rect 36452 17008 36504 17060
rect 38660 17051 38712 17060
rect 38660 17017 38669 17051
rect 38669 17017 38703 17051
rect 38703 17017 38712 17051
rect 38660 17008 38712 17017
rect 5711 16838 5763 16890
rect 5775 16838 5827 16890
rect 5839 16838 5891 16890
rect 5903 16838 5955 16890
rect 5967 16838 6019 16890
rect 15233 16838 15285 16890
rect 15297 16838 15349 16890
rect 15361 16838 15413 16890
rect 15425 16838 15477 16890
rect 15489 16838 15541 16890
rect 24755 16838 24807 16890
rect 24819 16838 24871 16890
rect 24883 16838 24935 16890
rect 24947 16838 24999 16890
rect 25011 16838 25063 16890
rect 34277 16838 34329 16890
rect 34341 16838 34393 16890
rect 34405 16838 34457 16890
rect 34469 16838 34521 16890
rect 34533 16838 34585 16890
rect 5356 16736 5408 16788
rect 5448 16736 5500 16788
rect 6000 16736 6052 16788
rect 12532 16736 12584 16788
rect 13820 16736 13872 16788
rect 17224 16736 17276 16788
rect 17960 16736 18012 16788
rect 18144 16736 18196 16788
rect 20996 16736 21048 16788
rect 22284 16736 22336 16788
rect 26608 16779 26660 16788
rect 26608 16745 26617 16779
rect 26617 16745 26651 16779
rect 26651 16745 26660 16779
rect 26608 16736 26660 16745
rect 15384 16668 15436 16720
rect 4620 16600 4672 16652
rect 4896 16643 4948 16652
rect 4896 16609 4905 16643
rect 4905 16609 4939 16643
rect 4939 16609 4948 16643
rect 4896 16600 4948 16609
rect 11796 16600 11848 16652
rect 12256 16600 12308 16652
rect 2044 16532 2096 16584
rect 3148 16532 3200 16584
rect 5632 16532 5684 16584
rect 7748 16532 7800 16584
rect 9312 16532 9364 16584
rect 13820 16600 13872 16652
rect 940 16464 992 16516
rect 12256 16464 12308 16516
rect 13636 16575 13688 16584
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 15936 16600 15988 16652
rect 12900 16464 12952 16516
rect 14556 16464 14608 16516
rect 15108 16532 15160 16584
rect 15660 16464 15712 16516
rect 17224 16575 17276 16584
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 17316 16575 17368 16584
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 17316 16532 17368 16541
rect 20996 16643 21048 16652
rect 20996 16609 21005 16643
rect 21005 16609 21039 16643
rect 21039 16609 21048 16643
rect 20996 16600 21048 16609
rect 23020 16600 23072 16652
rect 23572 16600 23624 16652
rect 25136 16668 25188 16720
rect 25320 16643 25372 16652
rect 25320 16609 25329 16643
rect 25329 16609 25363 16643
rect 25363 16609 25372 16643
rect 25320 16600 25372 16609
rect 25780 16600 25832 16652
rect 30656 16643 30708 16652
rect 30656 16609 30665 16643
rect 30665 16609 30699 16643
rect 30699 16609 30708 16643
rect 30656 16600 30708 16609
rect 32864 16668 32916 16720
rect 32680 16600 32732 16652
rect 35072 16600 35124 16652
rect 23848 16532 23900 16584
rect 26332 16532 26384 16584
rect 27344 16575 27396 16584
rect 27344 16541 27353 16575
rect 27353 16541 27387 16575
rect 27387 16541 27396 16575
rect 27344 16532 27396 16541
rect 28908 16532 28960 16584
rect 30840 16532 30892 16584
rect 2688 16439 2740 16448
rect 2688 16405 2697 16439
rect 2697 16405 2731 16439
rect 2731 16405 2740 16439
rect 2688 16396 2740 16405
rect 3240 16396 3292 16448
rect 4344 16439 4396 16448
rect 4344 16405 4353 16439
rect 4353 16405 4387 16439
rect 4387 16405 4396 16439
rect 4344 16396 4396 16405
rect 4436 16396 4488 16448
rect 4988 16396 5040 16448
rect 5448 16396 5500 16448
rect 12716 16396 12768 16448
rect 16028 16396 16080 16448
rect 16304 16507 16356 16516
rect 16304 16473 16313 16507
rect 16313 16473 16347 16507
rect 16347 16473 16356 16507
rect 16304 16464 16356 16473
rect 20720 16464 20772 16516
rect 22284 16464 22336 16516
rect 24492 16464 24544 16516
rect 16764 16396 16816 16448
rect 17960 16439 18012 16448
rect 17960 16405 17969 16439
rect 17969 16405 18003 16439
rect 18003 16405 18012 16439
rect 17960 16396 18012 16405
rect 22744 16439 22796 16448
rect 22744 16405 22753 16439
rect 22753 16405 22787 16439
rect 22787 16405 22796 16439
rect 22744 16396 22796 16405
rect 23204 16439 23256 16448
rect 23204 16405 23213 16439
rect 23213 16405 23247 16439
rect 23247 16405 23256 16439
rect 23204 16396 23256 16405
rect 23756 16396 23808 16448
rect 27620 16507 27672 16516
rect 27620 16473 27629 16507
rect 27629 16473 27663 16507
rect 27663 16473 27672 16507
rect 27620 16464 27672 16473
rect 32312 16464 32364 16516
rect 32956 16464 33008 16516
rect 33232 16575 33284 16584
rect 33232 16541 33241 16575
rect 33241 16541 33275 16575
rect 33275 16541 33284 16575
rect 33232 16532 33284 16541
rect 33508 16575 33560 16584
rect 33508 16541 33517 16575
rect 33517 16541 33551 16575
rect 33551 16541 33560 16575
rect 33508 16532 33560 16541
rect 33968 16532 34020 16584
rect 35256 16575 35308 16584
rect 35256 16541 35265 16575
rect 35265 16541 35299 16575
rect 35299 16541 35308 16575
rect 35256 16532 35308 16541
rect 35532 16532 35584 16584
rect 36636 16532 36688 16584
rect 34336 16464 34388 16516
rect 35164 16507 35216 16516
rect 35164 16473 35173 16507
rect 35173 16473 35207 16507
rect 35207 16473 35216 16507
rect 35164 16464 35216 16473
rect 25228 16396 25280 16448
rect 28908 16396 28960 16448
rect 29000 16396 29052 16448
rect 29920 16396 29972 16448
rect 30472 16396 30524 16448
rect 32772 16396 32824 16448
rect 33232 16396 33284 16448
rect 33692 16396 33744 16448
rect 33876 16396 33928 16448
rect 36360 16396 36412 16448
rect 10472 16294 10524 16346
rect 10536 16294 10588 16346
rect 10600 16294 10652 16346
rect 10664 16294 10716 16346
rect 10728 16294 10780 16346
rect 19994 16294 20046 16346
rect 20058 16294 20110 16346
rect 20122 16294 20174 16346
rect 20186 16294 20238 16346
rect 20250 16294 20302 16346
rect 29516 16294 29568 16346
rect 29580 16294 29632 16346
rect 29644 16294 29696 16346
rect 29708 16294 29760 16346
rect 29772 16294 29824 16346
rect 39038 16294 39090 16346
rect 39102 16294 39154 16346
rect 39166 16294 39218 16346
rect 39230 16294 39282 16346
rect 39294 16294 39346 16346
rect 2688 16192 2740 16244
rect 8576 16192 8628 16244
rect 3240 16124 3292 16176
rect 5632 16167 5684 16176
rect 5632 16133 5641 16167
rect 5641 16133 5675 16167
rect 5675 16133 5684 16167
rect 5632 16124 5684 16133
rect 6828 16124 6880 16176
rect 10968 16192 11020 16244
rect 9128 16167 9180 16176
rect 9128 16133 9137 16167
rect 9137 16133 9171 16167
rect 9171 16133 9180 16167
rect 9128 16124 9180 16133
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 4528 16056 4580 16108
rect 2228 16031 2280 16040
rect 2228 15997 2237 16031
rect 2237 15997 2271 16031
rect 2271 15997 2280 16031
rect 2228 15988 2280 15997
rect 2504 16031 2556 16040
rect 2504 15997 2513 16031
rect 2513 15997 2547 16031
rect 2547 15997 2556 16031
rect 2504 15988 2556 15997
rect 5172 15988 5224 16040
rect 7748 15988 7800 16040
rect 8668 15963 8720 15972
rect 8668 15929 8677 15963
rect 8677 15929 8711 15963
rect 8711 15929 8720 15963
rect 8668 15920 8720 15929
rect 9680 16056 9732 16108
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 11704 16192 11756 16244
rect 12716 16192 12768 16244
rect 21824 16192 21876 16244
rect 12624 16124 12676 16176
rect 13544 16167 13596 16176
rect 13544 16133 13553 16167
rect 13553 16133 13587 16167
rect 13587 16133 13596 16167
rect 13544 16124 13596 16133
rect 14188 16124 14240 16176
rect 15108 16124 15160 16176
rect 23204 16192 23256 16244
rect 23572 16192 23624 16244
rect 27528 16192 27580 16244
rect 29184 16235 29236 16244
rect 29184 16201 29193 16235
rect 29193 16201 29227 16235
rect 29227 16201 29236 16235
rect 29184 16192 29236 16201
rect 29920 16167 29972 16176
rect 29920 16133 29929 16167
rect 29929 16133 29963 16167
rect 29963 16133 29972 16167
rect 29920 16124 29972 16133
rect 30932 16124 30984 16176
rect 11796 16056 11848 16108
rect 13176 16056 13228 16108
rect 15384 16056 15436 16108
rect 16028 16099 16080 16108
rect 16028 16065 16037 16099
rect 16037 16065 16071 16099
rect 16071 16065 16080 16099
rect 16028 16056 16080 16065
rect 16396 16056 16448 16108
rect 20352 16056 20404 16108
rect 27344 16056 27396 16108
rect 2964 15852 3016 15904
rect 3148 15852 3200 15904
rect 10048 15852 10100 15904
rect 11060 15963 11112 15972
rect 11060 15929 11069 15963
rect 11069 15929 11103 15963
rect 11103 15929 11112 15963
rect 11060 15920 11112 15929
rect 11888 15852 11940 15904
rect 12716 15963 12768 15972
rect 12716 15929 12725 15963
rect 12725 15929 12759 15963
rect 12759 15929 12768 15963
rect 12716 15920 12768 15929
rect 12900 15920 12952 15972
rect 14004 15852 14056 15904
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 15752 15988 15804 16040
rect 16304 16031 16356 16040
rect 16304 15997 16313 16031
rect 16313 15997 16347 16031
rect 16347 15997 16356 16031
rect 16304 15988 16356 15997
rect 20720 15988 20772 16040
rect 22376 15988 22428 16040
rect 26700 15988 26752 16040
rect 29368 15988 29420 16040
rect 33692 16192 33744 16244
rect 35348 16192 35400 16244
rect 31300 16056 31352 16108
rect 33048 16124 33100 16176
rect 33324 16124 33376 16176
rect 34704 16124 34756 16176
rect 35072 16124 35124 16176
rect 38476 16124 38528 16176
rect 32956 16056 33008 16108
rect 35808 16099 35860 16108
rect 35808 16065 35817 16099
rect 35817 16065 35851 16099
rect 35851 16065 35860 16099
rect 35808 16056 35860 16065
rect 15200 15920 15252 15972
rect 17868 15920 17920 15972
rect 19892 15852 19944 15904
rect 22744 15852 22796 15904
rect 28724 15852 28776 15904
rect 33876 15988 33928 16040
rect 34152 15988 34204 16040
rect 36636 16099 36688 16108
rect 36636 16065 36645 16099
rect 36645 16065 36679 16099
rect 36679 16065 36688 16099
rect 36636 16056 36688 16065
rect 37188 16056 37240 16108
rect 37556 16056 37608 16108
rect 30932 15920 30984 15972
rect 30288 15852 30340 15904
rect 30656 15852 30708 15904
rect 32588 15895 32640 15904
rect 32588 15861 32597 15895
rect 32597 15861 32631 15895
rect 32631 15861 32640 15895
rect 32588 15852 32640 15861
rect 34796 15920 34848 15972
rect 37924 15988 37976 16040
rect 34152 15852 34204 15904
rect 34888 15895 34940 15904
rect 34888 15861 34897 15895
rect 34897 15861 34931 15895
rect 34931 15861 34940 15895
rect 34888 15852 34940 15861
rect 35440 15895 35492 15904
rect 35440 15861 35449 15895
rect 35449 15861 35483 15895
rect 35483 15861 35492 15895
rect 35440 15852 35492 15861
rect 36728 15895 36780 15904
rect 36728 15861 36737 15895
rect 36737 15861 36771 15895
rect 36771 15861 36780 15895
rect 36728 15852 36780 15861
rect 37280 15852 37332 15904
rect 5711 15750 5763 15802
rect 5775 15750 5827 15802
rect 5839 15750 5891 15802
rect 5903 15750 5955 15802
rect 5967 15750 6019 15802
rect 15233 15750 15285 15802
rect 15297 15750 15349 15802
rect 15361 15750 15413 15802
rect 15425 15750 15477 15802
rect 15489 15750 15541 15802
rect 24755 15750 24807 15802
rect 24819 15750 24871 15802
rect 24883 15750 24935 15802
rect 24947 15750 24999 15802
rect 25011 15750 25063 15802
rect 34277 15750 34329 15802
rect 34341 15750 34393 15802
rect 34405 15750 34457 15802
rect 34469 15750 34521 15802
rect 34533 15750 34585 15802
rect 2504 15648 2556 15700
rect 3608 15648 3660 15700
rect 3148 15555 3200 15564
rect 3148 15521 3157 15555
rect 3157 15521 3191 15555
rect 3191 15521 3200 15555
rect 3148 15512 3200 15521
rect 3332 15555 3384 15564
rect 3332 15521 3341 15555
rect 3341 15521 3375 15555
rect 3375 15521 3384 15555
rect 3332 15512 3384 15521
rect 4620 15512 4672 15564
rect 8208 15691 8260 15700
rect 8208 15657 8217 15691
rect 8217 15657 8251 15691
rect 8251 15657 8260 15691
rect 8208 15648 8260 15657
rect 11704 15648 11756 15700
rect 11888 15648 11940 15700
rect 13636 15648 13688 15700
rect 13728 15691 13780 15700
rect 13728 15657 13737 15691
rect 13737 15657 13771 15691
rect 13771 15657 13780 15691
rect 13728 15648 13780 15657
rect 14188 15648 14240 15700
rect 15108 15648 15160 15700
rect 9772 15555 9824 15564
rect 9772 15521 9781 15555
rect 9781 15521 9815 15555
rect 9815 15521 9824 15555
rect 9772 15512 9824 15521
rect 12624 15512 12676 15564
rect 12900 15512 12952 15564
rect 19984 15580 20036 15632
rect 20628 15580 20680 15632
rect 24860 15580 24912 15632
rect 26424 15691 26476 15700
rect 26424 15657 26433 15691
rect 26433 15657 26467 15691
rect 26467 15657 26476 15691
rect 26424 15648 26476 15657
rect 27620 15648 27672 15700
rect 28724 15648 28776 15700
rect 30932 15648 30984 15700
rect 31208 15648 31260 15700
rect 35992 15648 36044 15700
rect 14096 15512 14148 15564
rect 16856 15512 16908 15564
rect 940 15444 992 15496
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 5632 15444 5684 15496
rect 6644 15444 6696 15496
rect 7564 15444 7616 15496
rect 9680 15444 9732 15496
rect 14372 15444 14424 15496
rect 17960 15444 18012 15496
rect 2688 15376 2740 15428
rect 4160 15376 4212 15428
rect 4712 15376 4764 15428
rect 12348 15376 12400 15428
rect 14280 15419 14332 15428
rect 14280 15385 14289 15419
rect 14289 15385 14323 15419
rect 14323 15385 14332 15419
rect 14280 15376 14332 15385
rect 15016 15419 15068 15428
rect 3056 15351 3108 15360
rect 3056 15317 3065 15351
rect 3065 15317 3099 15351
rect 3099 15317 3108 15351
rect 3056 15308 3108 15317
rect 8208 15308 8260 15360
rect 8300 15308 8352 15360
rect 10140 15308 10192 15360
rect 11888 15308 11940 15360
rect 12624 15308 12676 15360
rect 15016 15385 15025 15419
rect 15025 15385 15059 15419
rect 15059 15385 15068 15419
rect 15016 15376 15068 15385
rect 20352 15444 20404 15496
rect 20720 15444 20772 15496
rect 23848 15487 23900 15496
rect 23848 15453 23857 15487
rect 23857 15453 23891 15487
rect 23891 15453 23900 15487
rect 23848 15444 23900 15453
rect 26608 15512 26660 15564
rect 26240 15444 26292 15496
rect 26332 15487 26384 15496
rect 26332 15453 26341 15487
rect 26341 15453 26375 15487
rect 26375 15453 26384 15487
rect 26332 15444 26384 15453
rect 28172 15580 28224 15632
rect 28540 15580 28592 15632
rect 28908 15555 28960 15564
rect 28908 15521 28917 15555
rect 28917 15521 28951 15555
rect 28951 15521 28960 15555
rect 28908 15512 28960 15521
rect 31300 15580 31352 15632
rect 31760 15580 31812 15632
rect 32956 15580 33008 15632
rect 30196 15555 30248 15564
rect 30196 15521 30205 15555
rect 30205 15521 30239 15555
rect 30239 15521 30248 15555
rect 30196 15512 30248 15521
rect 29920 15487 29972 15496
rect 29920 15453 29929 15487
rect 29929 15453 29963 15487
rect 29963 15453 29972 15487
rect 29920 15444 29972 15453
rect 31392 15487 31444 15496
rect 31392 15453 31401 15487
rect 31401 15453 31435 15487
rect 31435 15453 31444 15487
rect 31392 15444 31444 15453
rect 31484 15444 31536 15496
rect 14832 15308 14884 15360
rect 19156 15376 19208 15428
rect 19708 15376 19760 15428
rect 20076 15376 20128 15428
rect 20904 15376 20956 15428
rect 17684 15351 17736 15360
rect 17684 15317 17693 15351
rect 17693 15317 17727 15351
rect 17727 15317 17736 15351
rect 17684 15308 17736 15317
rect 17960 15308 18012 15360
rect 19432 15308 19484 15360
rect 21824 15376 21876 15428
rect 25504 15376 25556 15428
rect 25780 15419 25832 15428
rect 25780 15385 25789 15419
rect 25789 15385 25823 15419
rect 25823 15385 25832 15419
rect 25780 15376 25832 15385
rect 26700 15376 26752 15428
rect 31576 15419 31628 15428
rect 31576 15385 31585 15419
rect 31585 15385 31619 15419
rect 31619 15385 31628 15419
rect 31576 15376 31628 15385
rect 23940 15351 23992 15360
rect 23940 15317 23949 15351
rect 23949 15317 23983 15351
rect 23983 15317 23992 15351
rect 23940 15308 23992 15317
rect 25688 15351 25740 15360
rect 25688 15317 25697 15351
rect 25697 15317 25731 15351
rect 25731 15317 25740 15351
rect 25688 15308 25740 15317
rect 28816 15308 28868 15360
rect 31116 15308 31168 15360
rect 32220 15444 32272 15496
rect 33784 15512 33836 15564
rect 33232 15487 33284 15496
rect 33232 15453 33241 15487
rect 33241 15453 33275 15487
rect 33275 15453 33284 15487
rect 33232 15444 33284 15453
rect 33508 15444 33560 15496
rect 35072 15555 35124 15564
rect 35072 15521 35081 15555
rect 35081 15521 35115 15555
rect 35115 15521 35124 15555
rect 35072 15512 35124 15521
rect 36452 15580 36504 15632
rect 37372 15512 37424 15564
rect 37924 15487 37976 15496
rect 37924 15453 37933 15487
rect 37933 15453 37967 15487
rect 37967 15453 37976 15487
rect 37924 15444 37976 15453
rect 34152 15376 34204 15428
rect 32036 15308 32088 15360
rect 32128 15308 32180 15360
rect 33232 15308 33284 15360
rect 33416 15308 33468 15360
rect 36728 15376 36780 15428
rect 37096 15419 37148 15428
rect 37096 15385 37105 15419
rect 37105 15385 37139 15419
rect 37139 15385 37148 15419
rect 37096 15376 37148 15385
rect 10472 15206 10524 15258
rect 10536 15206 10588 15258
rect 10600 15206 10652 15258
rect 10664 15206 10716 15258
rect 10728 15206 10780 15258
rect 19994 15206 20046 15258
rect 20058 15206 20110 15258
rect 20122 15206 20174 15258
rect 20186 15206 20238 15258
rect 20250 15206 20302 15258
rect 29516 15206 29568 15258
rect 29580 15206 29632 15258
rect 29644 15206 29696 15258
rect 29708 15206 29760 15258
rect 29772 15206 29824 15258
rect 39038 15206 39090 15258
rect 39102 15206 39154 15258
rect 39166 15206 39218 15258
rect 39230 15206 39282 15258
rect 39294 15206 39346 15258
rect 4896 15104 4948 15156
rect 4988 15104 5040 15156
rect 2596 15036 2648 15088
rect 4252 15036 4304 15088
rect 5540 15079 5592 15088
rect 5540 15045 5549 15079
rect 5549 15045 5583 15079
rect 5583 15045 5592 15079
rect 5540 15036 5592 15045
rect 5632 15036 5684 15088
rect 6368 15036 6420 15088
rect 2320 14900 2372 14952
rect 2228 14832 2280 14884
rect 3976 14900 4028 14952
rect 5264 14875 5316 14884
rect 5264 14841 5273 14875
rect 5273 14841 5307 14875
rect 5307 14841 5316 14875
rect 5264 14832 5316 14841
rect 5356 14832 5408 14884
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 7932 15147 7984 15156
rect 7932 15113 7941 15147
rect 7941 15113 7975 15147
rect 7975 15113 7984 15147
rect 7932 15104 7984 15113
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 11244 15104 11296 15156
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 11888 15104 11940 15156
rect 12256 15104 12308 15156
rect 11152 15036 11204 15088
rect 11428 15036 11480 15088
rect 11980 15036 12032 15088
rect 18052 15104 18104 15156
rect 18236 15104 18288 15156
rect 18512 15147 18564 15156
rect 18512 15113 18521 15147
rect 18521 15113 18555 15147
rect 18555 15113 18564 15147
rect 18512 15104 18564 15113
rect 21088 15147 21140 15156
rect 21088 15113 21097 15147
rect 21097 15113 21131 15147
rect 21131 15113 21140 15147
rect 21088 15104 21140 15113
rect 8392 14968 8444 15020
rect 11796 14968 11848 15020
rect 12072 15011 12124 15020
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 8116 14900 8168 14952
rect 8300 14900 8352 14952
rect 9864 14900 9916 14952
rect 11520 14900 11572 14952
rect 12348 14900 12400 14952
rect 12716 14900 12768 14952
rect 14096 15079 14148 15088
rect 14096 15045 14105 15079
rect 14105 15045 14139 15079
rect 14139 15045 14148 15079
rect 14096 15036 14148 15045
rect 16672 15036 16724 15088
rect 17500 15036 17552 15088
rect 13728 14968 13780 15020
rect 14372 14900 14424 14952
rect 15844 14968 15896 15020
rect 19432 15036 19484 15088
rect 19984 15036 20036 15088
rect 16028 14900 16080 14952
rect 16396 14900 16448 14952
rect 17224 14900 17276 14952
rect 17500 14943 17552 14952
rect 17500 14909 17509 14943
rect 17509 14909 17543 14943
rect 17543 14909 17552 14943
rect 17500 14900 17552 14909
rect 18604 14900 18656 14952
rect 1952 14764 2004 14816
rect 3056 14764 3108 14816
rect 5540 14764 5592 14816
rect 6276 14764 6328 14816
rect 13544 14832 13596 14884
rect 16948 14875 17000 14884
rect 16948 14841 16957 14875
rect 16957 14841 16991 14875
rect 16991 14841 17000 14875
rect 16948 14832 17000 14841
rect 17868 14832 17920 14884
rect 19432 14900 19484 14952
rect 20628 14968 20680 15020
rect 21364 14943 21416 14952
rect 21364 14909 21373 14943
rect 21373 14909 21407 14943
rect 21407 14909 21416 14943
rect 21364 14900 21416 14909
rect 22928 15104 22980 15156
rect 31668 15104 31720 15156
rect 22192 15036 22244 15088
rect 23296 15036 23348 15088
rect 23940 15036 23992 15088
rect 26240 15036 26292 15088
rect 31392 15036 31444 15088
rect 22100 14900 22152 14952
rect 26792 14968 26844 15020
rect 28264 15011 28316 15020
rect 28264 14977 28273 15011
rect 28273 14977 28307 15011
rect 28307 14977 28316 15011
rect 28264 14968 28316 14977
rect 28448 15011 28500 15020
rect 28448 14977 28457 15011
rect 28457 14977 28491 15011
rect 28491 14977 28500 15011
rect 28448 14968 28500 14977
rect 28540 15011 28592 15020
rect 28540 14977 28549 15011
rect 28549 14977 28583 15011
rect 28583 14977 28592 15011
rect 28540 14968 28592 14977
rect 20628 14832 20680 14884
rect 25136 14943 25188 14952
rect 25136 14909 25145 14943
rect 25145 14909 25179 14943
rect 25179 14909 25188 14943
rect 25136 14900 25188 14909
rect 28356 14900 28408 14952
rect 28816 14968 28868 15020
rect 29092 14968 29144 15020
rect 32680 15104 32732 15156
rect 32864 15104 32916 15156
rect 32588 15036 32640 15088
rect 35072 15036 35124 15088
rect 35164 15079 35216 15088
rect 35164 15045 35173 15079
rect 35173 15045 35207 15079
rect 35207 15045 35216 15079
rect 35164 15036 35216 15045
rect 35900 15036 35952 15088
rect 38476 15079 38528 15088
rect 38476 15045 38485 15079
rect 38485 15045 38519 15079
rect 38519 15045 38528 15079
rect 38476 15036 38528 15045
rect 32312 15011 32364 15020
rect 32312 14977 32321 15011
rect 32321 14977 32355 15011
rect 32355 14977 32364 15011
rect 32312 14968 32364 14977
rect 34888 15011 34940 15020
rect 34888 14977 34897 15011
rect 34897 14977 34931 15011
rect 34931 14977 34940 15011
rect 34888 14968 34940 14977
rect 37832 14968 37884 15020
rect 38660 15011 38712 15020
rect 38660 14977 38669 15011
rect 38669 14977 38703 15011
rect 38703 14977 38712 15011
rect 38660 14968 38712 14977
rect 29920 14943 29972 14952
rect 29920 14909 29929 14943
rect 29929 14909 29963 14943
rect 29963 14909 29972 14943
rect 29920 14900 29972 14909
rect 30288 14900 30340 14952
rect 31024 14900 31076 14952
rect 32588 14943 32640 14952
rect 32588 14909 32597 14943
rect 32597 14909 32631 14943
rect 32631 14909 32640 14943
rect 32588 14900 32640 14909
rect 32680 14900 32732 14952
rect 33968 14900 34020 14952
rect 11244 14764 11296 14816
rect 11612 14764 11664 14816
rect 13084 14764 13136 14816
rect 18420 14764 18472 14816
rect 21088 14764 21140 14816
rect 26332 14764 26384 14816
rect 28448 14764 28500 14816
rect 31116 14764 31168 14816
rect 31760 14764 31812 14816
rect 36636 14807 36688 14816
rect 36636 14773 36645 14807
rect 36645 14773 36679 14807
rect 36679 14773 36688 14807
rect 36636 14764 36688 14773
rect 5711 14662 5763 14714
rect 5775 14662 5827 14714
rect 5839 14662 5891 14714
rect 5903 14662 5955 14714
rect 5967 14662 6019 14714
rect 15233 14662 15285 14714
rect 15297 14662 15349 14714
rect 15361 14662 15413 14714
rect 15425 14662 15477 14714
rect 15489 14662 15541 14714
rect 24755 14662 24807 14714
rect 24819 14662 24871 14714
rect 24883 14662 24935 14714
rect 24947 14662 24999 14714
rect 25011 14662 25063 14714
rect 34277 14662 34329 14714
rect 34341 14662 34393 14714
rect 34405 14662 34457 14714
rect 34469 14662 34521 14714
rect 34533 14662 34585 14714
rect 1768 14603 1820 14612
rect 1768 14569 1777 14603
rect 1777 14569 1811 14603
rect 1811 14569 1820 14603
rect 1768 14560 1820 14569
rect 2136 14603 2188 14612
rect 2136 14569 2145 14603
rect 2145 14569 2179 14603
rect 2179 14569 2188 14603
rect 2136 14560 2188 14569
rect 2596 14560 2648 14612
rect 4988 14560 5040 14612
rect 6736 14560 6788 14612
rect 8760 14560 8812 14612
rect 2320 14424 2372 14476
rect 3056 14424 3108 14476
rect 9220 14492 9272 14544
rect 3976 14424 4028 14476
rect 7012 14424 7064 14476
rect 9956 14492 10008 14544
rect 1676 14331 1728 14340
rect 1676 14297 1685 14331
rect 1685 14297 1719 14331
rect 1719 14297 1728 14331
rect 1676 14288 1728 14297
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 3700 14356 3752 14408
rect 4344 14356 4396 14408
rect 9588 14467 9640 14476
rect 9588 14433 9597 14467
rect 9597 14433 9631 14467
rect 9631 14433 9640 14467
rect 9588 14424 9640 14433
rect 13268 14492 13320 14544
rect 13452 14492 13504 14544
rect 14556 14560 14608 14612
rect 10876 14467 10928 14476
rect 10876 14433 10885 14467
rect 10885 14433 10919 14467
rect 10919 14433 10928 14467
rect 10876 14424 10928 14433
rect 7196 14399 7248 14408
rect 7196 14365 7205 14399
rect 7205 14365 7239 14399
rect 7239 14365 7248 14399
rect 12716 14424 12768 14476
rect 7196 14356 7248 14365
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 11888 14356 11940 14408
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 13268 14399 13320 14408
rect 13268 14365 13275 14399
rect 13275 14365 13320 14399
rect 13268 14356 13320 14365
rect 13912 14356 13964 14408
rect 14096 14356 14148 14408
rect 14464 14356 14516 14408
rect 14832 14399 14884 14408
rect 14832 14365 14841 14399
rect 14841 14365 14875 14399
rect 14875 14365 14884 14399
rect 14832 14356 14884 14365
rect 15016 14356 15068 14408
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 17500 14560 17552 14612
rect 17868 14560 17920 14612
rect 18788 14492 18840 14544
rect 17868 14424 17920 14476
rect 22100 14492 22152 14544
rect 26792 14560 26844 14612
rect 27804 14492 27856 14544
rect 27988 14492 28040 14544
rect 32312 14492 32364 14544
rect 34888 14492 34940 14544
rect 3148 14288 3200 14340
rect 3608 14288 3660 14340
rect 5172 14288 5224 14340
rect 6552 14288 6604 14340
rect 6644 14220 6696 14272
rect 6736 14263 6788 14272
rect 6736 14229 6745 14263
rect 6745 14229 6779 14263
rect 6779 14229 6788 14263
rect 6736 14220 6788 14229
rect 7104 14220 7156 14272
rect 8944 14288 8996 14340
rect 12072 14288 12124 14340
rect 12256 14331 12308 14340
rect 12256 14297 12265 14331
rect 12265 14297 12299 14331
rect 12299 14297 12308 14331
rect 12256 14288 12308 14297
rect 12992 14288 13044 14340
rect 13452 14331 13504 14340
rect 13452 14297 13461 14331
rect 13461 14297 13495 14331
rect 13495 14297 13504 14331
rect 13452 14288 13504 14297
rect 15660 14288 15712 14340
rect 16212 14288 16264 14340
rect 16672 14288 16724 14340
rect 8576 14220 8628 14272
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 17592 14288 17644 14340
rect 18512 14288 18564 14340
rect 20628 14424 20680 14476
rect 24860 14424 24912 14476
rect 25320 14424 25372 14476
rect 27620 14424 27672 14476
rect 28908 14467 28960 14476
rect 28908 14433 28917 14467
rect 28917 14433 28951 14467
rect 28951 14433 28960 14467
rect 28908 14424 28960 14433
rect 29000 14467 29052 14476
rect 29000 14433 29009 14467
rect 29009 14433 29043 14467
rect 29043 14433 29052 14467
rect 29000 14424 29052 14433
rect 29276 14424 29328 14476
rect 30472 14424 30524 14476
rect 31024 14467 31076 14476
rect 31024 14433 31033 14467
rect 31033 14433 31067 14467
rect 31067 14433 31076 14467
rect 31024 14424 31076 14433
rect 37372 14535 37424 14544
rect 37372 14501 37381 14535
rect 37381 14501 37415 14535
rect 37415 14501 37424 14535
rect 37372 14492 37424 14501
rect 19892 14356 19944 14408
rect 20720 14356 20772 14408
rect 30196 14356 30248 14408
rect 33140 14356 33192 14408
rect 33508 14356 33560 14408
rect 36360 14356 36412 14408
rect 37188 14399 37240 14408
rect 37188 14365 37197 14399
rect 37197 14365 37231 14399
rect 37231 14365 37240 14399
rect 37188 14356 37240 14365
rect 38108 14356 38160 14408
rect 21088 14331 21140 14340
rect 21088 14297 21097 14331
rect 21097 14297 21131 14331
rect 21131 14297 21140 14331
rect 21088 14288 21140 14297
rect 21180 14288 21232 14340
rect 23664 14288 23716 14340
rect 23848 14220 23900 14272
rect 28724 14288 28776 14340
rect 29920 14288 29972 14340
rect 30748 14288 30800 14340
rect 31300 14331 31352 14340
rect 31300 14297 31309 14331
rect 31309 14297 31343 14331
rect 31343 14297 31352 14331
rect 31300 14288 31352 14297
rect 26700 14220 26752 14272
rect 26792 14263 26844 14272
rect 26792 14229 26801 14263
rect 26801 14229 26835 14263
rect 26835 14229 26844 14263
rect 26792 14220 26844 14229
rect 28448 14263 28500 14272
rect 28448 14229 28457 14263
rect 28457 14229 28491 14263
rect 28491 14229 28500 14263
rect 28448 14220 28500 14229
rect 29000 14220 29052 14272
rect 29276 14220 29328 14272
rect 30012 14220 30064 14272
rect 31484 14220 31536 14272
rect 31576 14220 31628 14272
rect 35256 14331 35308 14340
rect 35256 14297 35265 14331
rect 35265 14297 35299 14331
rect 35299 14297 35308 14331
rect 35256 14288 35308 14297
rect 36636 14220 36688 14272
rect 36728 14263 36780 14272
rect 36728 14229 36737 14263
rect 36737 14229 36771 14263
rect 36771 14229 36780 14263
rect 36728 14220 36780 14229
rect 10472 14118 10524 14170
rect 10536 14118 10588 14170
rect 10600 14118 10652 14170
rect 10664 14118 10716 14170
rect 10728 14118 10780 14170
rect 19994 14118 20046 14170
rect 20058 14118 20110 14170
rect 20122 14118 20174 14170
rect 20186 14118 20238 14170
rect 20250 14118 20302 14170
rect 29516 14118 29568 14170
rect 29580 14118 29632 14170
rect 29644 14118 29696 14170
rect 29708 14118 29760 14170
rect 29772 14118 29824 14170
rect 39038 14118 39090 14170
rect 39102 14118 39154 14170
rect 39166 14118 39218 14170
rect 39230 14118 39282 14170
rect 39294 14118 39346 14170
rect 2044 13991 2096 14000
rect 2044 13957 2053 13991
rect 2053 13957 2087 13991
rect 2087 13957 2096 13991
rect 2044 13948 2096 13957
rect 3424 13948 3476 14000
rect 6552 14016 6604 14068
rect 6644 14016 6696 14068
rect 8484 14016 8536 14068
rect 11612 14016 11664 14068
rect 3976 13880 4028 13932
rect 10048 13948 10100 14000
rect 14556 14016 14608 14068
rect 14372 13948 14424 14000
rect 14464 13948 14516 14000
rect 15016 14016 15068 14068
rect 15108 13948 15160 14000
rect 15568 13948 15620 14000
rect 16672 13948 16724 14000
rect 17592 13948 17644 14000
rect 5448 13880 5500 13932
rect 2136 13812 2188 13864
rect 3700 13812 3752 13864
rect 5540 13812 5592 13864
rect 4068 13676 4120 13728
rect 5632 13676 5684 13728
rect 6644 13676 6696 13728
rect 8024 13880 8076 13932
rect 8944 13880 8996 13932
rect 10508 13880 10560 13932
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 12624 13880 12676 13932
rect 7012 13812 7064 13864
rect 8300 13812 8352 13864
rect 8208 13744 8260 13796
rect 13452 13812 13504 13864
rect 14648 13880 14700 13932
rect 14832 13812 14884 13864
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 7196 13676 7248 13728
rect 8024 13676 8076 13728
rect 10324 13744 10376 13796
rect 10508 13744 10560 13796
rect 12532 13744 12584 13796
rect 12072 13719 12124 13728
rect 12072 13685 12081 13719
rect 12081 13685 12115 13719
rect 12115 13685 12124 13719
rect 12072 13676 12124 13685
rect 14648 13676 14700 13728
rect 15108 13676 15160 13728
rect 15660 13676 15712 13728
rect 16396 13880 16448 13932
rect 16672 13812 16724 13864
rect 18236 13880 18288 13932
rect 19708 13991 19760 14000
rect 19708 13957 19717 13991
rect 19717 13957 19751 13991
rect 19751 13957 19760 13991
rect 19708 13948 19760 13957
rect 20720 13948 20772 14000
rect 21088 13948 21140 14000
rect 25228 14016 25280 14068
rect 23480 13948 23532 14000
rect 23848 13948 23900 14000
rect 27896 14016 27948 14068
rect 17224 13744 17276 13796
rect 17408 13855 17460 13864
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 16672 13676 16724 13728
rect 16856 13719 16908 13728
rect 16856 13685 16865 13719
rect 16865 13685 16899 13719
rect 16899 13685 16908 13719
rect 16856 13676 16908 13685
rect 18236 13744 18288 13796
rect 20444 13880 20496 13932
rect 20628 13812 20680 13864
rect 18788 13744 18840 13796
rect 19432 13744 19484 13796
rect 21364 13880 21416 13932
rect 21640 13880 21692 13932
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 24860 13880 24912 13889
rect 27436 13880 27488 13932
rect 17684 13676 17736 13728
rect 17776 13676 17828 13728
rect 25136 13812 25188 13864
rect 27252 13855 27304 13864
rect 27252 13821 27261 13855
rect 27261 13821 27295 13855
rect 27295 13821 27304 13855
rect 27252 13812 27304 13821
rect 29368 14016 29420 14068
rect 29920 14059 29972 14068
rect 29920 14025 29929 14059
rect 29929 14025 29963 14059
rect 29963 14025 29972 14059
rect 29920 14016 29972 14025
rect 30380 14016 30432 14068
rect 30840 14016 30892 14068
rect 32680 14016 32732 14068
rect 33692 14016 33744 14068
rect 34612 14016 34664 14068
rect 34704 14059 34756 14068
rect 34704 14025 34713 14059
rect 34713 14025 34747 14059
rect 34747 14025 34756 14059
rect 34704 14016 34756 14025
rect 35256 14016 35308 14068
rect 28448 13991 28500 14000
rect 28448 13957 28457 13991
rect 28457 13957 28491 13991
rect 28491 13957 28500 13991
rect 28448 13948 28500 13957
rect 28724 13948 28776 14000
rect 30196 13880 30248 13932
rect 33324 13948 33376 14000
rect 34244 13948 34296 14000
rect 36728 14016 36780 14068
rect 36636 13948 36688 14000
rect 33048 13880 33100 13932
rect 33692 13880 33744 13932
rect 21824 13744 21876 13796
rect 21088 13676 21140 13728
rect 22192 13676 22244 13728
rect 22468 13719 22520 13728
rect 22468 13685 22498 13719
rect 22498 13685 22520 13719
rect 22468 13676 22520 13685
rect 25872 13676 25924 13728
rect 26516 13676 26568 13728
rect 28080 13676 28132 13728
rect 28908 13676 28960 13728
rect 31852 13812 31904 13864
rect 32772 13855 32824 13864
rect 32772 13821 32781 13855
rect 32781 13821 32815 13855
rect 32815 13821 32824 13855
rect 32772 13812 32824 13821
rect 33140 13812 33192 13864
rect 33508 13812 33560 13864
rect 33968 13923 34020 13932
rect 33968 13889 33977 13923
rect 33977 13889 34011 13923
rect 34011 13889 34020 13923
rect 33968 13880 34020 13889
rect 35072 13880 35124 13932
rect 35900 13855 35952 13864
rect 35900 13821 35909 13855
rect 35909 13821 35943 13855
rect 35943 13821 35952 13855
rect 35900 13812 35952 13821
rect 34244 13744 34296 13796
rect 35716 13744 35768 13796
rect 36820 13855 36872 13864
rect 36820 13821 36829 13855
rect 36829 13821 36863 13855
rect 36863 13821 36872 13855
rect 36820 13812 36872 13821
rect 38108 13923 38160 13932
rect 38108 13889 38117 13923
rect 38117 13889 38151 13923
rect 38151 13889 38160 13923
rect 38108 13880 38160 13889
rect 37832 13812 37884 13864
rect 36452 13744 36504 13796
rect 37280 13744 37332 13796
rect 33048 13676 33100 13728
rect 35624 13676 35676 13728
rect 38200 13719 38252 13728
rect 38200 13685 38209 13719
rect 38209 13685 38243 13719
rect 38243 13685 38252 13719
rect 38200 13676 38252 13685
rect 5711 13574 5763 13626
rect 5775 13574 5827 13626
rect 5839 13574 5891 13626
rect 5903 13574 5955 13626
rect 5967 13574 6019 13626
rect 15233 13574 15285 13626
rect 15297 13574 15349 13626
rect 15361 13574 15413 13626
rect 15425 13574 15477 13626
rect 15489 13574 15541 13626
rect 24755 13574 24807 13626
rect 24819 13574 24871 13626
rect 24883 13574 24935 13626
rect 24947 13574 24999 13626
rect 25011 13574 25063 13626
rect 34277 13574 34329 13626
rect 34341 13574 34393 13626
rect 34405 13574 34457 13626
rect 34469 13574 34521 13626
rect 34533 13574 34585 13626
rect 4068 13472 4120 13524
rect 2136 13404 2188 13456
rect 3700 13404 3752 13456
rect 1584 13268 1636 13320
rect 2044 13268 2096 13320
rect 3332 13311 3384 13320
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 5448 13336 5500 13388
rect 6552 13336 6604 13388
rect 6920 13336 6972 13388
rect 7288 13472 7340 13524
rect 8024 13472 8076 13524
rect 7472 13404 7524 13456
rect 14280 13472 14332 13524
rect 14556 13472 14608 13524
rect 14740 13515 14792 13524
rect 14740 13481 14749 13515
rect 14749 13481 14783 13515
rect 14783 13481 14792 13515
rect 14740 13472 14792 13481
rect 16120 13472 16172 13524
rect 16212 13472 16264 13524
rect 17132 13472 17184 13524
rect 17408 13472 17460 13524
rect 17776 13472 17828 13524
rect 18420 13515 18472 13524
rect 18420 13481 18429 13515
rect 18429 13481 18463 13515
rect 18463 13481 18472 13515
rect 18420 13472 18472 13481
rect 18788 13515 18840 13524
rect 18788 13481 18797 13515
rect 18797 13481 18831 13515
rect 18831 13481 18840 13515
rect 18788 13472 18840 13481
rect 21088 13472 21140 13524
rect 7748 13336 7800 13388
rect 9772 13336 9824 13388
rect 16580 13404 16632 13456
rect 19800 13404 19852 13456
rect 21824 13472 21876 13524
rect 22836 13472 22888 13524
rect 23020 13472 23072 13524
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 9864 13268 9916 13320
rect 12348 13336 12400 13388
rect 13268 13336 13320 13388
rect 13360 13336 13412 13388
rect 5356 13200 5408 13252
rect 6184 13243 6236 13252
rect 6184 13209 6193 13243
rect 6193 13209 6227 13243
rect 6227 13209 6236 13243
rect 6184 13200 6236 13209
rect 7840 13200 7892 13252
rect 940 13132 992 13184
rect 2504 13132 2556 13184
rect 4436 13175 4488 13184
rect 4436 13141 4445 13175
rect 4445 13141 4479 13175
rect 4479 13141 4488 13175
rect 4436 13132 4488 13141
rect 4620 13132 4672 13184
rect 6000 13132 6052 13184
rect 6368 13132 6420 13184
rect 8024 13132 8076 13184
rect 9956 13200 10008 13252
rect 8300 13175 8352 13184
rect 8300 13141 8325 13175
rect 8325 13141 8352 13175
rect 8300 13132 8352 13141
rect 8760 13132 8812 13184
rect 10876 13132 10928 13184
rect 11060 13243 11112 13252
rect 11060 13209 11069 13243
rect 11069 13209 11103 13243
rect 11103 13209 11112 13243
rect 11060 13200 11112 13209
rect 12072 13200 12124 13252
rect 13176 13311 13228 13320
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 13636 13268 13688 13320
rect 14924 13268 14976 13320
rect 15200 13336 15252 13388
rect 16028 13336 16080 13388
rect 16672 13336 16724 13388
rect 16856 13336 16908 13388
rect 15752 13268 15804 13320
rect 16120 13268 16172 13320
rect 12348 13132 12400 13184
rect 12440 13132 12492 13184
rect 13268 13200 13320 13252
rect 14280 13200 14332 13252
rect 15660 13200 15712 13252
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 18696 13268 18748 13320
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 19524 13268 19576 13320
rect 20720 13336 20772 13388
rect 21272 13336 21324 13388
rect 27436 13404 27488 13456
rect 26148 13336 26200 13388
rect 26608 13379 26660 13388
rect 26608 13345 26617 13379
rect 26617 13345 26651 13379
rect 26651 13345 26660 13379
rect 26608 13336 26660 13345
rect 27712 13336 27764 13388
rect 27988 13379 28040 13388
rect 27988 13345 27997 13379
rect 27997 13345 28031 13379
rect 28031 13345 28040 13379
rect 27988 13336 28040 13345
rect 22192 13268 22244 13320
rect 22376 13268 22428 13320
rect 22744 13268 22796 13320
rect 22836 13268 22888 13320
rect 16948 13200 17000 13252
rect 17684 13200 17736 13252
rect 18144 13243 18196 13252
rect 18144 13209 18153 13243
rect 18153 13209 18187 13243
rect 18187 13209 18196 13243
rect 18144 13200 18196 13209
rect 18236 13200 18288 13252
rect 18420 13200 18472 13252
rect 20444 13200 20496 13252
rect 14740 13132 14792 13184
rect 14924 13132 14976 13184
rect 15292 13132 15344 13184
rect 16764 13132 16816 13184
rect 19892 13132 19944 13184
rect 20352 13132 20404 13184
rect 22008 13200 22060 13252
rect 22560 13200 22612 13252
rect 23296 13200 23348 13252
rect 23848 13311 23900 13320
rect 23848 13277 23857 13311
rect 23857 13277 23891 13311
rect 23891 13277 23900 13311
rect 23848 13268 23900 13277
rect 24584 13268 24636 13320
rect 28908 13404 28960 13456
rect 30288 13404 30340 13456
rect 32772 13472 32824 13524
rect 33048 13472 33100 13524
rect 33692 13472 33744 13524
rect 33968 13404 34020 13456
rect 34060 13447 34112 13456
rect 34060 13413 34069 13447
rect 34069 13413 34103 13447
rect 34103 13413 34112 13447
rect 34060 13404 34112 13413
rect 29920 13336 29972 13388
rect 30932 13336 30984 13388
rect 32404 13336 32456 13388
rect 34796 13336 34848 13388
rect 34888 13379 34940 13388
rect 34888 13345 34897 13379
rect 34897 13345 34931 13379
rect 34931 13345 34940 13379
rect 34888 13336 34940 13345
rect 22192 13132 22244 13184
rect 23664 13132 23716 13184
rect 23940 13175 23992 13184
rect 23940 13141 23949 13175
rect 23949 13141 23983 13175
rect 23983 13141 23992 13175
rect 23940 13132 23992 13141
rect 25596 13200 25648 13252
rect 30196 13268 30248 13320
rect 33692 13268 33744 13320
rect 33876 13268 33928 13320
rect 38384 13268 38436 13320
rect 26792 13200 26844 13252
rect 28172 13200 28224 13252
rect 30840 13243 30892 13252
rect 30840 13209 30849 13243
rect 30849 13209 30883 13243
rect 30883 13209 30892 13243
rect 30840 13200 30892 13209
rect 31852 13200 31904 13252
rect 25872 13132 25924 13184
rect 26516 13175 26568 13184
rect 26516 13141 26525 13175
rect 26525 13141 26559 13175
rect 26559 13141 26568 13175
rect 26516 13132 26568 13141
rect 28448 13132 28500 13184
rect 28816 13132 28868 13184
rect 30472 13132 30524 13184
rect 38200 13200 38252 13252
rect 39396 13200 39448 13252
rect 32864 13132 32916 13184
rect 35900 13132 35952 13184
rect 37372 13132 37424 13184
rect 37740 13132 37792 13184
rect 10472 13030 10524 13082
rect 10536 13030 10588 13082
rect 10600 13030 10652 13082
rect 10664 13030 10716 13082
rect 10728 13030 10780 13082
rect 19994 13030 20046 13082
rect 20058 13030 20110 13082
rect 20122 13030 20174 13082
rect 20186 13030 20238 13082
rect 20250 13030 20302 13082
rect 29516 13030 29568 13082
rect 29580 13030 29632 13082
rect 29644 13030 29696 13082
rect 29708 13030 29760 13082
rect 29772 13030 29824 13082
rect 39038 13030 39090 13082
rect 39102 13030 39154 13082
rect 39166 13030 39218 13082
rect 39230 13030 39282 13082
rect 39294 13030 39346 13082
rect 6092 12928 6144 12980
rect 6184 12928 6236 12980
rect 7748 12928 7800 12980
rect 8024 12971 8076 12980
rect 8024 12937 8033 12971
rect 8033 12937 8067 12971
rect 8067 12937 8076 12971
rect 8024 12928 8076 12937
rect 8300 12928 8352 12980
rect 3516 12860 3568 12912
rect 3792 12860 3844 12912
rect 4436 12860 4488 12912
rect 2044 12792 2096 12844
rect 5172 12835 5224 12844
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 1952 12656 2004 12708
rect 4528 12724 4580 12776
rect 3608 12656 3660 12708
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5632 12792 5684 12844
rect 7564 12792 7616 12844
rect 7840 12860 7892 12912
rect 11060 12928 11112 12980
rect 13176 12903 13228 12912
rect 13176 12869 13185 12903
rect 13185 12869 13219 12903
rect 13219 12869 13228 12903
rect 13176 12860 13228 12869
rect 13268 12860 13320 12912
rect 13544 12971 13596 12980
rect 13544 12937 13553 12971
rect 13553 12937 13587 12971
rect 13587 12937 13596 12971
rect 13544 12928 13596 12937
rect 14648 12928 14700 12980
rect 14924 12928 14976 12980
rect 15200 12928 15252 12980
rect 16396 12928 16448 12980
rect 16488 12928 16540 12980
rect 16764 12928 16816 12980
rect 18696 12928 18748 12980
rect 18880 12928 18932 12980
rect 7196 12656 7248 12708
rect 7472 12724 7524 12776
rect 8208 12767 8260 12776
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 9680 12835 9732 12844
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 9956 12792 10008 12844
rect 10140 12792 10192 12844
rect 10508 12792 10560 12844
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 12164 12835 12216 12844
rect 12164 12801 12173 12835
rect 12173 12801 12207 12835
rect 12207 12801 12216 12835
rect 12164 12792 12216 12801
rect 12900 12792 12952 12844
rect 13820 12792 13872 12844
rect 15108 12792 15160 12844
rect 15660 12792 15712 12844
rect 15844 12792 15896 12844
rect 10876 12724 10928 12776
rect 13728 12724 13780 12776
rect 15752 12724 15804 12776
rect 15936 12724 15988 12776
rect 18972 12860 19024 12912
rect 20720 12928 20772 12980
rect 25504 12928 25556 12980
rect 26240 12928 26292 12980
rect 26516 12928 26568 12980
rect 21272 12792 21324 12844
rect 21916 12792 21968 12844
rect 22836 12860 22888 12912
rect 23112 12860 23164 12912
rect 26148 12860 26200 12912
rect 27988 12903 28040 12912
rect 27988 12869 27997 12903
rect 27997 12869 28031 12903
rect 28031 12869 28040 12903
rect 27988 12860 28040 12869
rect 28356 12860 28408 12912
rect 31484 12971 31536 12980
rect 31484 12937 31493 12971
rect 31493 12937 31527 12971
rect 31527 12937 31536 12971
rect 31484 12928 31536 12937
rect 31760 12928 31812 12980
rect 32864 12928 32916 12980
rect 33140 12928 33192 12980
rect 33416 12928 33468 12980
rect 22376 12792 22428 12844
rect 22928 12835 22980 12844
rect 22928 12801 22937 12835
rect 22937 12801 22971 12835
rect 22971 12801 22980 12835
rect 22928 12792 22980 12801
rect 24492 12792 24544 12844
rect 25872 12792 25924 12844
rect 26240 12835 26292 12844
rect 26240 12801 26249 12835
rect 26249 12801 26283 12835
rect 26283 12801 26292 12835
rect 26240 12792 26292 12801
rect 28080 12792 28132 12844
rect 28264 12792 28316 12844
rect 28724 12835 28776 12844
rect 28724 12801 28733 12835
rect 28733 12801 28767 12835
rect 28767 12801 28776 12835
rect 28724 12792 28776 12801
rect 29092 12835 29144 12844
rect 29092 12801 29101 12835
rect 29101 12801 29135 12835
rect 29135 12801 29144 12835
rect 29092 12792 29144 12801
rect 29368 12792 29420 12844
rect 29920 12860 29972 12912
rect 30012 12903 30064 12912
rect 30012 12869 30021 12903
rect 30021 12869 30055 12903
rect 30055 12869 30064 12903
rect 30012 12860 30064 12869
rect 32680 12860 32732 12912
rect 35256 12928 35308 12980
rect 35440 12928 35492 12980
rect 22192 12767 22244 12776
rect 22192 12733 22201 12767
rect 22201 12733 22235 12767
rect 22235 12733 22244 12767
rect 22192 12724 22244 12733
rect 26608 12724 26660 12776
rect 28816 12724 28868 12776
rect 5264 12631 5316 12640
rect 5264 12597 5273 12631
rect 5273 12597 5307 12631
rect 5307 12597 5316 12631
rect 5264 12588 5316 12597
rect 9220 12588 9272 12640
rect 9680 12656 9732 12708
rect 10140 12588 10192 12640
rect 11520 12656 11572 12708
rect 12256 12656 12308 12708
rect 14648 12656 14700 12708
rect 10784 12588 10836 12640
rect 12348 12588 12400 12640
rect 12532 12588 12584 12640
rect 15476 12588 15528 12640
rect 22376 12656 22428 12708
rect 24216 12656 24268 12708
rect 31760 12724 31812 12776
rect 33048 12835 33100 12844
rect 33048 12801 33057 12835
rect 33057 12801 33091 12835
rect 33091 12801 33100 12835
rect 33048 12792 33100 12801
rect 35624 12860 35676 12912
rect 33324 12792 33376 12844
rect 33968 12792 34020 12844
rect 32864 12724 32916 12776
rect 35256 12792 35308 12844
rect 37464 12792 37516 12844
rect 37832 12792 37884 12844
rect 34888 12724 34940 12776
rect 16580 12588 16632 12640
rect 16948 12588 17000 12640
rect 17776 12588 17828 12640
rect 18328 12588 18380 12640
rect 18604 12588 18656 12640
rect 20444 12588 20496 12640
rect 25504 12588 25556 12640
rect 25688 12588 25740 12640
rect 25872 12588 25924 12640
rect 27436 12588 27488 12640
rect 30748 12588 30800 12640
rect 33324 12631 33376 12640
rect 33324 12597 33333 12631
rect 33333 12597 33367 12631
rect 33367 12597 33376 12631
rect 33324 12588 33376 12597
rect 33876 12631 33928 12640
rect 33876 12597 33885 12631
rect 33885 12597 33919 12631
rect 33919 12597 33928 12631
rect 33876 12588 33928 12597
rect 34152 12588 34204 12640
rect 34888 12588 34940 12640
rect 35256 12588 35308 12640
rect 38292 12631 38344 12640
rect 38292 12597 38301 12631
rect 38301 12597 38335 12631
rect 38335 12597 38344 12631
rect 38292 12588 38344 12597
rect 5711 12486 5763 12538
rect 5775 12486 5827 12538
rect 5839 12486 5891 12538
rect 5903 12486 5955 12538
rect 5967 12486 6019 12538
rect 15233 12486 15285 12538
rect 15297 12486 15349 12538
rect 15361 12486 15413 12538
rect 15425 12486 15477 12538
rect 15489 12486 15541 12538
rect 24755 12486 24807 12538
rect 24819 12486 24871 12538
rect 24883 12486 24935 12538
rect 24947 12486 24999 12538
rect 25011 12486 25063 12538
rect 34277 12486 34329 12538
rect 34341 12486 34393 12538
rect 34405 12486 34457 12538
rect 34469 12486 34521 12538
rect 34533 12486 34585 12538
rect 1768 12384 1820 12436
rect 3608 12384 3660 12436
rect 9956 12384 10008 12436
rect 10232 12384 10284 12436
rect 10600 12384 10652 12436
rect 2044 12248 2096 12300
rect 3148 12248 3200 12300
rect 5816 12248 5868 12300
rect 7012 12248 7064 12300
rect 8944 12316 8996 12368
rect 9128 12316 9180 12368
rect 10784 12316 10836 12368
rect 11244 12316 11296 12368
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 15568 12384 15620 12436
rect 16396 12384 16448 12436
rect 17776 12427 17828 12436
rect 17776 12393 17785 12427
rect 17785 12393 17819 12427
rect 17819 12393 17828 12427
rect 17776 12384 17828 12393
rect 20352 12427 20404 12436
rect 20352 12393 20361 12427
rect 20361 12393 20395 12427
rect 20395 12393 20404 12427
rect 20352 12384 20404 12393
rect 21088 12384 21140 12436
rect 21272 12427 21324 12436
rect 21272 12393 21281 12427
rect 21281 12393 21315 12427
rect 21315 12393 21324 12427
rect 21272 12384 21324 12393
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 5632 12180 5684 12232
rect 2688 12087 2740 12096
rect 2688 12053 2697 12087
rect 2697 12053 2731 12087
rect 2731 12053 2740 12087
rect 2688 12044 2740 12053
rect 3240 12044 3292 12096
rect 3884 12112 3936 12164
rect 7380 12155 7432 12164
rect 7380 12121 7389 12155
rect 7389 12121 7423 12155
rect 7423 12121 7432 12155
rect 7380 12112 7432 12121
rect 7748 12180 7800 12232
rect 8944 12180 8996 12232
rect 7840 12112 7892 12164
rect 6184 12044 6236 12096
rect 6460 12044 6512 12096
rect 9404 12112 9456 12164
rect 9864 12180 9916 12232
rect 10508 12180 10560 12232
rect 11244 12180 11296 12232
rect 11428 12180 11480 12232
rect 11888 12180 11940 12232
rect 9956 12112 10008 12164
rect 8668 12044 8720 12096
rect 9680 12044 9732 12096
rect 10600 12112 10652 12164
rect 17224 12316 17276 12368
rect 17316 12316 17368 12368
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 14004 12180 14056 12232
rect 14740 12180 14792 12232
rect 14832 12180 14884 12232
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 16488 12291 16540 12300
rect 16488 12257 16497 12291
rect 16497 12257 16531 12291
rect 16531 12257 16540 12291
rect 16488 12248 16540 12257
rect 16764 12248 16816 12300
rect 17408 12248 17460 12300
rect 17684 12316 17736 12368
rect 17960 12316 18012 12368
rect 19708 12316 19760 12368
rect 18696 12248 18748 12300
rect 19340 12248 19392 12300
rect 23112 12384 23164 12436
rect 23664 12384 23716 12436
rect 26056 12384 26108 12436
rect 26700 12384 26752 12436
rect 27436 12384 27488 12436
rect 21456 12316 21508 12368
rect 21640 12316 21692 12368
rect 10232 12044 10284 12096
rect 10784 12044 10836 12096
rect 11152 12044 11204 12096
rect 11612 12087 11664 12096
rect 11612 12053 11621 12087
rect 11621 12053 11655 12087
rect 11655 12053 11664 12087
rect 11612 12044 11664 12053
rect 11704 12044 11756 12096
rect 13268 12112 13320 12164
rect 13636 12112 13688 12164
rect 13728 12112 13780 12164
rect 16212 12112 16264 12164
rect 17684 12180 17736 12232
rect 17868 12112 17920 12164
rect 13912 12044 13964 12096
rect 14740 12044 14792 12096
rect 16028 12044 16080 12096
rect 16764 12044 16816 12096
rect 18420 12044 18472 12096
rect 20536 12180 20588 12232
rect 20720 12180 20772 12232
rect 25136 12248 25188 12300
rect 25964 12248 26016 12300
rect 21640 12180 21692 12232
rect 22652 12180 22704 12232
rect 23204 12180 23256 12232
rect 23848 12223 23900 12232
rect 23848 12189 23857 12223
rect 23857 12189 23891 12223
rect 23891 12189 23900 12223
rect 23848 12180 23900 12189
rect 24492 12180 24544 12232
rect 24584 12180 24636 12232
rect 27344 12180 27396 12232
rect 27896 12180 27948 12232
rect 29000 12384 29052 12436
rect 31116 12384 31168 12436
rect 33048 12384 33100 12436
rect 34888 12384 34940 12436
rect 35072 12427 35124 12436
rect 35072 12393 35081 12427
rect 35081 12393 35115 12427
rect 35115 12393 35124 12427
rect 35072 12384 35124 12393
rect 35992 12427 36044 12436
rect 35992 12393 36001 12427
rect 36001 12393 36035 12427
rect 36035 12393 36044 12427
rect 35992 12384 36044 12393
rect 37188 12384 37240 12436
rect 31668 12316 31720 12368
rect 33140 12316 33192 12368
rect 28356 12248 28408 12300
rect 28632 12248 28684 12300
rect 29368 12248 29420 12300
rect 31760 12248 31812 12300
rect 32864 12248 32916 12300
rect 33416 12248 33468 12300
rect 33692 12248 33744 12300
rect 35072 12248 35124 12300
rect 20812 12112 20864 12164
rect 20996 12112 21048 12164
rect 21548 12112 21600 12164
rect 22560 12112 22612 12164
rect 23020 12112 23072 12164
rect 25412 12112 25464 12164
rect 20628 12044 20680 12096
rect 21088 12044 21140 12096
rect 21456 12044 21508 12096
rect 21824 12044 21876 12096
rect 24492 12044 24544 12096
rect 25688 12044 25740 12096
rect 27252 12112 27304 12164
rect 29276 12112 29328 12164
rect 30012 12112 30064 12164
rect 26976 12044 27028 12096
rect 27344 12044 27396 12096
rect 27528 12044 27580 12096
rect 28724 12044 28776 12096
rect 28908 12044 28960 12096
rect 29920 12044 29972 12096
rect 30380 12044 30432 12096
rect 30564 12044 30616 12096
rect 31392 12044 31444 12096
rect 31484 12044 31536 12096
rect 32312 12044 32364 12096
rect 32772 12112 32824 12164
rect 33048 12112 33100 12164
rect 33140 12112 33192 12164
rect 34152 12112 34204 12164
rect 32588 12087 32640 12096
rect 32588 12053 32613 12087
rect 32613 12053 32640 12087
rect 32588 12044 32640 12053
rect 32864 12044 32916 12096
rect 34612 12180 34664 12232
rect 35900 12223 35952 12232
rect 35900 12189 35909 12223
rect 35909 12189 35943 12223
rect 35943 12189 35952 12223
rect 35900 12180 35952 12189
rect 37464 12248 37516 12300
rect 38016 12180 38068 12232
rect 38384 12180 38436 12232
rect 34796 12112 34848 12164
rect 35164 12112 35216 12164
rect 36084 12044 36136 12096
rect 36820 12044 36872 12096
rect 10472 11942 10524 11994
rect 10536 11942 10588 11994
rect 10600 11942 10652 11994
rect 10664 11942 10716 11994
rect 10728 11942 10780 11994
rect 19994 11942 20046 11994
rect 20058 11942 20110 11994
rect 20122 11942 20174 11994
rect 20186 11942 20238 11994
rect 20250 11942 20302 11994
rect 29516 11942 29568 11994
rect 29580 11942 29632 11994
rect 29644 11942 29696 11994
rect 29708 11942 29760 11994
rect 29772 11942 29824 11994
rect 39038 11942 39090 11994
rect 39102 11942 39154 11994
rect 39166 11942 39218 11994
rect 39230 11942 39282 11994
rect 39294 11942 39346 11994
rect 2228 11840 2280 11892
rect 1768 11747 1820 11756
rect 1768 11713 1777 11747
rect 1777 11713 1811 11747
rect 1811 11713 1820 11747
rect 1768 11704 1820 11713
rect 2872 11840 2924 11892
rect 3424 11840 3476 11892
rect 5356 11840 5408 11892
rect 5448 11840 5500 11892
rect 6644 11840 6696 11892
rect 7840 11840 7892 11892
rect 3792 11704 3844 11756
rect 6460 11772 6512 11824
rect 6828 11772 6880 11824
rect 9312 11840 9364 11892
rect 9772 11840 9824 11892
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 5540 11636 5592 11688
rect 7012 11704 7064 11756
rect 7288 11747 7340 11756
rect 7288 11713 7297 11747
rect 7297 11713 7331 11747
rect 7331 11713 7340 11747
rect 7288 11704 7340 11713
rect 7932 11704 7984 11756
rect 8300 11747 8352 11756
rect 8300 11713 8309 11747
rect 8309 11713 8343 11747
rect 8343 11713 8352 11747
rect 8300 11704 8352 11713
rect 5816 11679 5868 11688
rect 5816 11645 5825 11679
rect 5825 11645 5859 11679
rect 5859 11645 5868 11679
rect 5816 11636 5868 11645
rect 7380 11636 7432 11688
rect 8116 11636 8168 11688
rect 9864 11704 9916 11756
rect 10784 11704 10836 11756
rect 7748 11568 7800 11620
rect 8484 11568 8536 11620
rect 9588 11568 9640 11620
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 2044 11500 2096 11552
rect 2688 11500 2740 11552
rect 4252 11500 4304 11552
rect 6276 11500 6328 11552
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 9404 11500 9456 11552
rect 10324 11679 10376 11688
rect 10324 11645 10333 11679
rect 10333 11645 10367 11679
rect 10367 11645 10376 11679
rect 10324 11636 10376 11645
rect 10968 11840 11020 11892
rect 11244 11704 11296 11756
rect 13820 11840 13872 11892
rect 13912 11840 13964 11892
rect 15660 11840 15712 11892
rect 16856 11840 16908 11892
rect 13176 11815 13228 11824
rect 13176 11781 13185 11815
rect 13185 11781 13219 11815
rect 13219 11781 13228 11815
rect 13176 11772 13228 11781
rect 15844 11772 15896 11824
rect 12624 11704 12676 11756
rect 16028 11704 16080 11756
rect 17960 11840 18012 11892
rect 18696 11840 18748 11892
rect 18972 11840 19024 11892
rect 17500 11815 17552 11824
rect 17500 11781 17509 11815
rect 17509 11781 17543 11815
rect 17543 11781 17552 11815
rect 17500 11772 17552 11781
rect 18512 11772 18564 11824
rect 20444 11883 20496 11892
rect 20444 11849 20453 11883
rect 20453 11849 20487 11883
rect 20487 11849 20496 11883
rect 20444 11840 20496 11849
rect 20536 11883 20588 11892
rect 20536 11849 20545 11883
rect 20545 11849 20579 11883
rect 20579 11849 20588 11883
rect 20536 11840 20588 11849
rect 22376 11840 22428 11892
rect 17040 11704 17092 11756
rect 10416 11568 10468 11620
rect 12440 11568 12492 11620
rect 16212 11636 16264 11688
rect 16304 11636 16356 11688
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 17868 11704 17920 11756
rect 17960 11704 18012 11756
rect 18236 11704 18288 11756
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 19524 11704 19576 11756
rect 20444 11704 20496 11756
rect 21824 11772 21876 11824
rect 22100 11772 22152 11824
rect 22928 11772 22980 11824
rect 25136 11840 25188 11892
rect 21640 11704 21692 11756
rect 21732 11704 21784 11756
rect 19708 11636 19760 11688
rect 22652 11704 22704 11756
rect 23940 11772 23992 11824
rect 24768 11772 24820 11824
rect 26056 11840 26108 11892
rect 25780 11772 25832 11824
rect 26424 11772 26476 11824
rect 27528 11772 27580 11824
rect 28172 11772 28224 11824
rect 22468 11636 22520 11688
rect 25964 11704 26016 11756
rect 28908 11883 28960 11892
rect 28908 11849 28917 11883
rect 28917 11849 28951 11883
rect 28951 11849 28960 11883
rect 28908 11840 28960 11849
rect 29184 11840 29236 11892
rect 29460 11815 29512 11824
rect 29460 11781 29469 11815
rect 29469 11781 29503 11815
rect 29503 11781 29512 11815
rect 29460 11772 29512 11781
rect 30012 11772 30064 11824
rect 31760 11772 31812 11824
rect 32312 11772 32364 11824
rect 33416 11840 33468 11892
rect 30564 11704 30616 11756
rect 30748 11704 30800 11756
rect 31392 11704 31444 11756
rect 10876 11500 10928 11552
rect 12256 11500 12308 11552
rect 12992 11500 13044 11552
rect 13728 11500 13780 11552
rect 14464 11500 14516 11552
rect 15660 11500 15712 11552
rect 16672 11500 16724 11552
rect 18236 11543 18288 11552
rect 18236 11509 18245 11543
rect 18245 11509 18279 11543
rect 18279 11509 18288 11543
rect 18236 11500 18288 11509
rect 18420 11500 18472 11552
rect 20720 11500 20772 11552
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 21364 11500 21416 11509
rect 22376 11568 22428 11620
rect 22560 11543 22612 11552
rect 22560 11509 22569 11543
rect 22569 11509 22603 11543
rect 22603 11509 22612 11543
rect 22560 11500 22612 11509
rect 25596 11568 25648 11620
rect 26148 11636 26200 11688
rect 27896 11636 27948 11688
rect 29092 11636 29144 11688
rect 31116 11636 31168 11688
rect 31208 11679 31260 11688
rect 31208 11645 31217 11679
rect 31217 11645 31251 11679
rect 31251 11645 31260 11679
rect 31208 11636 31260 11645
rect 32128 11636 32180 11688
rect 32404 11704 32456 11756
rect 33048 11704 33100 11756
rect 32588 11636 32640 11688
rect 33140 11679 33192 11688
rect 33140 11645 33149 11679
rect 33149 11645 33183 11679
rect 33183 11645 33192 11679
rect 33140 11636 33192 11645
rect 33968 11704 34020 11756
rect 34796 11704 34848 11756
rect 38016 11747 38068 11756
rect 38016 11713 38025 11747
rect 38025 11713 38059 11747
rect 38059 11713 38068 11747
rect 38016 11704 38068 11713
rect 34612 11636 34664 11688
rect 26240 11568 26292 11620
rect 26884 11568 26936 11620
rect 28724 11568 28776 11620
rect 33324 11568 33376 11620
rect 35900 11636 35952 11688
rect 25136 11500 25188 11552
rect 25688 11500 25740 11552
rect 29368 11500 29420 11552
rect 29644 11543 29696 11552
rect 29644 11509 29653 11543
rect 29653 11509 29687 11543
rect 29687 11509 29696 11543
rect 29644 11500 29696 11509
rect 30564 11500 30616 11552
rect 33968 11543 34020 11552
rect 33968 11509 33977 11543
rect 33977 11509 34011 11543
rect 34011 11509 34020 11543
rect 33968 11500 34020 11509
rect 5711 11398 5763 11450
rect 5775 11398 5827 11450
rect 5839 11398 5891 11450
rect 5903 11398 5955 11450
rect 5967 11398 6019 11450
rect 15233 11398 15285 11450
rect 15297 11398 15349 11450
rect 15361 11398 15413 11450
rect 15425 11398 15477 11450
rect 15489 11398 15541 11450
rect 24755 11398 24807 11450
rect 24819 11398 24871 11450
rect 24883 11398 24935 11450
rect 24947 11398 24999 11450
rect 25011 11398 25063 11450
rect 34277 11398 34329 11450
rect 34341 11398 34393 11450
rect 34405 11398 34457 11450
rect 34469 11398 34521 11450
rect 34533 11398 34585 11450
rect 3884 11296 3936 11348
rect 4344 11296 4396 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 3056 11228 3108 11280
rect 3148 11203 3200 11212
rect 3148 11169 3157 11203
rect 3157 11169 3191 11203
rect 3191 11169 3200 11203
rect 3148 11160 3200 11169
rect 3424 11160 3476 11212
rect 5356 11228 5408 11280
rect 5632 11160 5684 11212
rect 940 11024 992 11076
rect 2872 11092 2924 11144
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 6000 11228 6052 11280
rect 6276 11228 6328 11280
rect 8116 11228 8168 11280
rect 8300 11228 8352 11280
rect 9128 11296 9180 11348
rect 10508 11296 10560 11348
rect 11612 11296 11664 11348
rect 12440 11296 12492 11348
rect 15660 11296 15712 11348
rect 16304 11296 16356 11348
rect 17132 11296 17184 11348
rect 17316 11296 17368 11348
rect 17500 11296 17552 11348
rect 13636 11228 13688 11280
rect 7656 11160 7708 11212
rect 9404 11203 9456 11212
rect 9404 11169 9413 11203
rect 9413 11169 9447 11203
rect 9447 11169 9456 11203
rect 9404 11160 9456 11169
rect 11888 11203 11940 11212
rect 11888 11169 11897 11203
rect 11897 11169 11931 11203
rect 11931 11169 11940 11203
rect 11888 11160 11940 11169
rect 12624 11160 12676 11212
rect 18236 11228 18288 11280
rect 18420 11296 18472 11348
rect 19616 11296 19668 11348
rect 16028 11160 16080 11212
rect 17408 11160 17460 11212
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 6828 11092 6880 11144
rect 7472 11092 7524 11144
rect 7748 11135 7800 11144
rect 7748 11101 7757 11135
rect 7757 11101 7791 11135
rect 7791 11101 7800 11135
rect 7748 11092 7800 11101
rect 8484 11092 8536 11144
rect 8944 11092 8996 11144
rect 11796 11092 11848 11144
rect 11980 11092 12032 11144
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 17960 11092 18012 11144
rect 21640 11296 21692 11348
rect 21824 11296 21876 11348
rect 22652 11296 22704 11348
rect 23940 11339 23992 11348
rect 23940 11305 23949 11339
rect 23949 11305 23983 11339
rect 23983 11305 23992 11339
rect 23940 11296 23992 11305
rect 20720 11203 20772 11212
rect 20720 11169 20729 11203
rect 20729 11169 20763 11203
rect 20763 11169 20772 11203
rect 20720 11160 20772 11169
rect 25136 11228 25188 11280
rect 25596 11296 25648 11348
rect 26332 11296 26384 11348
rect 20536 11135 20588 11144
rect 20536 11101 20545 11135
rect 20545 11101 20579 11135
rect 20579 11101 20588 11135
rect 20536 11092 20588 11101
rect 23756 11092 23808 11144
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 23848 11092 23900 11101
rect 24584 11092 24636 11144
rect 25688 11228 25740 11280
rect 26056 11160 26108 11212
rect 26424 11160 26476 11212
rect 3884 11024 3936 11076
rect 4252 11067 4304 11076
rect 4252 11033 4261 11067
rect 4261 11033 4295 11067
rect 4295 11033 4304 11067
rect 4252 11024 4304 11033
rect 5632 11024 5684 11076
rect 6092 10956 6144 11008
rect 6828 10956 6880 11008
rect 9312 10956 9364 11008
rect 10232 10956 10284 11008
rect 11888 10956 11940 11008
rect 16212 11024 16264 11076
rect 18512 11024 18564 11076
rect 23020 11067 23072 11076
rect 23020 11033 23029 11067
rect 23029 11033 23063 11067
rect 23063 11033 23072 11067
rect 23020 11024 23072 11033
rect 23572 11024 23624 11076
rect 24308 11024 24360 11076
rect 26240 11092 26292 11144
rect 26608 11296 26660 11348
rect 28264 11296 28316 11348
rect 29276 11296 29328 11348
rect 29460 11296 29512 11348
rect 31300 11296 31352 11348
rect 34980 11339 35032 11348
rect 34980 11305 34989 11339
rect 34989 11305 35023 11339
rect 35023 11305 35032 11339
rect 34980 11296 35032 11305
rect 36084 11296 36136 11348
rect 27160 11228 27212 11280
rect 27528 11228 27580 11280
rect 28816 11228 28868 11280
rect 32036 11271 32088 11280
rect 32036 11237 32045 11271
rect 32045 11237 32079 11271
rect 32079 11237 32088 11271
rect 32036 11228 32088 11237
rect 32404 11228 32456 11280
rect 32588 11228 32640 11280
rect 34152 11228 34204 11280
rect 35992 11228 36044 11280
rect 26608 11160 26660 11212
rect 27896 11203 27948 11212
rect 27896 11169 27905 11203
rect 27905 11169 27939 11203
rect 27939 11169 27948 11203
rect 27896 11160 27948 11169
rect 30380 11160 30432 11212
rect 31208 11203 31260 11212
rect 31208 11169 31217 11203
rect 31217 11169 31251 11203
rect 31251 11169 31260 11203
rect 31208 11160 31260 11169
rect 31760 11160 31812 11212
rect 26884 11092 26936 11144
rect 28540 11092 28592 11144
rect 28724 11092 28776 11144
rect 30012 11092 30064 11144
rect 30196 11092 30248 11144
rect 32588 11135 32640 11144
rect 32588 11101 32597 11135
rect 32597 11101 32631 11135
rect 32631 11101 32640 11135
rect 32588 11092 32640 11101
rect 36268 11160 36320 11212
rect 37464 11092 37516 11144
rect 38108 11092 38160 11144
rect 16764 10999 16816 11008
rect 16764 10965 16773 10999
rect 16773 10965 16807 10999
rect 16807 10965 16816 10999
rect 16764 10956 16816 10965
rect 17132 10999 17184 11008
rect 17132 10965 17141 10999
rect 17141 10965 17175 10999
rect 17175 10965 17184 10999
rect 17132 10956 17184 10965
rect 19432 10956 19484 11008
rect 21732 10956 21784 11008
rect 24216 10956 24268 11008
rect 26424 11024 26476 11076
rect 25596 10999 25648 11008
rect 25596 10965 25605 10999
rect 25605 10965 25639 10999
rect 25639 10965 25648 10999
rect 25596 10956 25648 10965
rect 25780 10956 25832 11008
rect 26792 11024 26844 11076
rect 27712 11024 27764 11076
rect 26884 10999 26936 11008
rect 26884 10965 26893 10999
rect 26893 10965 26927 10999
rect 26927 10965 26936 10999
rect 26884 10956 26936 10965
rect 27160 10956 27212 11008
rect 28172 10999 28224 11008
rect 28172 10965 28181 10999
rect 28181 10965 28215 10999
rect 28215 10965 28224 10999
rect 28172 10956 28224 10965
rect 29184 11024 29236 11076
rect 29644 11024 29696 11076
rect 31024 11024 31076 11076
rect 31300 11024 31352 11076
rect 31576 11024 31628 11076
rect 32864 11067 32916 11076
rect 32864 11033 32873 11067
rect 32873 11033 32907 11067
rect 32907 11033 32916 11067
rect 32864 11024 32916 11033
rect 33876 11024 33928 11076
rect 34428 11024 34480 11076
rect 30564 10956 30616 11008
rect 31484 10956 31536 11008
rect 32128 10956 32180 11008
rect 36452 10956 36504 11008
rect 37648 11067 37700 11076
rect 37648 11033 37657 11067
rect 37657 11033 37691 11067
rect 37691 11033 37700 11067
rect 37648 11024 37700 11033
rect 39396 11024 39448 11076
rect 37740 10956 37792 11008
rect 10472 10854 10524 10906
rect 10536 10854 10588 10906
rect 10600 10854 10652 10906
rect 10664 10854 10716 10906
rect 10728 10854 10780 10906
rect 19994 10854 20046 10906
rect 20058 10854 20110 10906
rect 20122 10854 20174 10906
rect 20186 10854 20238 10906
rect 20250 10854 20302 10906
rect 29516 10854 29568 10906
rect 29580 10854 29632 10906
rect 29644 10854 29696 10906
rect 29708 10854 29760 10906
rect 29772 10854 29824 10906
rect 39038 10854 39090 10906
rect 39102 10854 39154 10906
rect 39166 10854 39218 10906
rect 39230 10854 39282 10906
rect 39294 10854 39346 10906
rect 5264 10752 5316 10804
rect 5356 10752 5408 10804
rect 8208 10752 8260 10804
rect 8852 10752 8904 10804
rect 1952 10684 2004 10736
rect 2412 10684 2464 10736
rect 5724 10684 5776 10736
rect 6736 10684 6788 10736
rect 8024 10684 8076 10736
rect 9404 10752 9456 10804
rect 10048 10684 10100 10736
rect 2872 10659 2924 10668
rect 2872 10625 2881 10659
rect 2881 10625 2915 10659
rect 2915 10625 2924 10659
rect 2872 10616 2924 10625
rect 6920 10616 6972 10668
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 9036 10616 9088 10668
rect 9404 10616 9456 10668
rect 10232 10616 10284 10668
rect 11060 10616 11112 10668
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 12072 10684 12124 10736
rect 13452 10684 13504 10736
rect 14464 10795 14516 10804
rect 14464 10761 14473 10795
rect 14473 10761 14507 10795
rect 14507 10761 14516 10795
rect 14464 10752 14516 10761
rect 14924 10752 14976 10804
rect 15384 10795 15436 10804
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 15568 10752 15620 10804
rect 16672 10684 16724 10736
rect 18604 10752 18656 10804
rect 22284 10752 22336 10804
rect 17500 10684 17552 10736
rect 21364 10684 21416 10736
rect 2320 10548 2372 10600
rect 3884 10548 3936 10600
rect 3792 10412 3844 10464
rect 6000 10523 6052 10532
rect 6000 10489 6009 10523
rect 6009 10489 6043 10523
rect 6043 10489 6052 10523
rect 6000 10480 6052 10489
rect 8944 10480 8996 10532
rect 12624 10548 12676 10600
rect 9128 10480 9180 10532
rect 10232 10480 10284 10532
rect 7104 10412 7156 10464
rect 11428 10412 11480 10464
rect 12072 10455 12124 10464
rect 12072 10421 12081 10455
rect 12081 10421 12115 10455
rect 12115 10421 12124 10455
rect 12072 10412 12124 10421
rect 13452 10548 13504 10600
rect 14464 10548 14516 10600
rect 16488 10548 16540 10600
rect 17316 10548 17368 10600
rect 17408 10591 17460 10600
rect 17408 10557 17417 10591
rect 17417 10557 17451 10591
rect 17451 10557 17460 10591
rect 17408 10548 17460 10557
rect 17500 10480 17552 10532
rect 13728 10412 13780 10464
rect 17132 10412 17184 10464
rect 19800 10616 19852 10668
rect 20628 10616 20680 10668
rect 23848 10752 23900 10804
rect 23940 10752 23992 10804
rect 24768 10684 24820 10736
rect 25964 10752 26016 10804
rect 25596 10616 25648 10668
rect 28172 10684 28224 10736
rect 29276 10752 29328 10804
rect 32680 10752 32732 10804
rect 33600 10752 33652 10804
rect 33876 10752 33928 10804
rect 34980 10752 35032 10804
rect 35716 10752 35768 10804
rect 29552 10684 29604 10736
rect 32312 10684 32364 10736
rect 34428 10684 34480 10736
rect 37372 10684 37424 10736
rect 17868 10548 17920 10600
rect 21272 10548 21324 10600
rect 20628 10480 20680 10532
rect 24492 10548 24544 10600
rect 25044 10548 25096 10600
rect 25136 10548 25188 10600
rect 26240 10659 26292 10668
rect 26240 10625 26249 10659
rect 26249 10625 26283 10659
rect 26283 10625 26292 10659
rect 26240 10616 26292 10625
rect 26332 10659 26384 10668
rect 26332 10625 26341 10659
rect 26341 10625 26375 10659
rect 26375 10625 26384 10659
rect 26332 10616 26384 10625
rect 27068 10616 27120 10668
rect 27436 10616 27488 10668
rect 28264 10616 28316 10668
rect 30564 10616 30616 10668
rect 31392 10659 31444 10668
rect 31392 10625 31401 10659
rect 31401 10625 31435 10659
rect 31435 10625 31444 10659
rect 31392 10616 31444 10625
rect 18788 10412 18840 10464
rect 24400 10480 24452 10532
rect 26700 10548 26752 10600
rect 27252 10548 27304 10600
rect 27160 10480 27212 10532
rect 23664 10412 23716 10464
rect 25504 10412 25556 10464
rect 25596 10412 25648 10464
rect 26240 10412 26292 10464
rect 28080 10412 28132 10464
rect 29092 10548 29144 10600
rect 31852 10616 31904 10668
rect 34520 10659 34572 10668
rect 34520 10625 34529 10659
rect 34529 10625 34563 10659
rect 34563 10625 34572 10659
rect 34520 10616 34572 10625
rect 37832 10616 37884 10668
rect 38016 10616 38068 10668
rect 38384 10616 38436 10668
rect 30472 10480 30524 10532
rect 31208 10480 31260 10532
rect 32588 10548 32640 10600
rect 34796 10591 34848 10600
rect 34796 10557 34805 10591
rect 34805 10557 34839 10591
rect 34839 10557 34848 10591
rect 34796 10548 34848 10557
rect 33692 10480 33744 10532
rect 34152 10480 34204 10532
rect 30196 10412 30248 10464
rect 31392 10412 31444 10464
rect 32128 10412 32180 10464
rect 33600 10412 33652 10464
rect 35808 10412 35860 10464
rect 36636 10412 36688 10464
rect 37648 10412 37700 10464
rect 38200 10455 38252 10464
rect 38200 10421 38209 10455
rect 38209 10421 38243 10455
rect 38243 10421 38252 10455
rect 38200 10412 38252 10421
rect 5711 10310 5763 10362
rect 5775 10310 5827 10362
rect 5839 10310 5891 10362
rect 5903 10310 5955 10362
rect 5967 10310 6019 10362
rect 15233 10310 15285 10362
rect 15297 10310 15349 10362
rect 15361 10310 15413 10362
rect 15425 10310 15477 10362
rect 15489 10310 15541 10362
rect 24755 10310 24807 10362
rect 24819 10310 24871 10362
rect 24883 10310 24935 10362
rect 24947 10310 24999 10362
rect 25011 10310 25063 10362
rect 34277 10310 34329 10362
rect 34341 10310 34393 10362
rect 34405 10310 34457 10362
rect 34469 10310 34521 10362
rect 34533 10310 34585 10362
rect 2688 10208 2740 10260
rect 5356 10208 5408 10260
rect 5632 10251 5684 10260
rect 5632 10217 5641 10251
rect 5641 10217 5675 10251
rect 5675 10217 5684 10251
rect 5632 10208 5684 10217
rect 8944 10208 8996 10260
rect 9680 10208 9732 10260
rect 10048 10208 10100 10260
rect 10232 10208 10284 10260
rect 1768 10004 1820 10056
rect 2596 10072 2648 10124
rect 4896 10072 4948 10124
rect 5816 10072 5868 10124
rect 6552 10072 6604 10124
rect 9312 10140 9364 10192
rect 11060 10140 11112 10192
rect 14096 10208 14148 10260
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 8852 10072 8904 10124
rect 5172 10004 5224 10056
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 6276 10004 6328 10056
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 8208 10004 8260 10056
rect 9312 10004 9364 10056
rect 11336 10004 11388 10056
rect 12900 10140 12952 10192
rect 13084 10140 13136 10192
rect 12808 10072 12860 10124
rect 16488 10140 16540 10192
rect 16764 10140 16816 10192
rect 18512 10251 18564 10260
rect 18512 10217 18521 10251
rect 18521 10217 18555 10251
rect 18555 10217 18564 10251
rect 18512 10208 18564 10217
rect 20720 10208 20772 10260
rect 14924 10072 14976 10124
rect 2228 9979 2280 9988
rect 2228 9945 2237 9979
rect 2237 9945 2271 9979
rect 2271 9945 2280 9979
rect 2228 9936 2280 9945
rect 2596 9979 2648 9988
rect 2596 9945 2605 9979
rect 2605 9945 2639 9979
rect 2639 9945 2648 9979
rect 2596 9936 2648 9945
rect 4436 9936 4488 9988
rect 6092 9936 6144 9988
rect 7104 9979 7156 9988
rect 7104 9945 7113 9979
rect 7113 9945 7147 9979
rect 7147 9945 7156 9979
rect 7104 9936 7156 9945
rect 9864 9979 9916 9988
rect 9864 9945 9873 9979
rect 9873 9945 9907 9979
rect 9907 9945 9916 9979
rect 9864 9936 9916 9945
rect 11152 9936 11204 9988
rect 11888 9936 11940 9988
rect 13452 9936 13504 9988
rect 13544 9936 13596 9988
rect 14832 10004 14884 10056
rect 17408 10072 17460 10124
rect 17684 10072 17736 10124
rect 19708 10072 19760 10124
rect 20628 10115 20680 10124
rect 20628 10081 20637 10115
rect 20637 10081 20671 10115
rect 20671 10081 20680 10115
rect 20628 10072 20680 10081
rect 21640 10072 21692 10124
rect 16304 10004 16356 10056
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 19340 10004 19392 10056
rect 15660 9936 15712 9988
rect 16212 9936 16264 9988
rect 1032 9868 1084 9920
rect 4160 9911 4212 9920
rect 4160 9877 4169 9911
rect 4169 9877 4203 9911
rect 4203 9877 4212 9911
rect 4160 9868 4212 9877
rect 4528 9911 4580 9920
rect 4528 9877 4537 9911
rect 4537 9877 4571 9911
rect 4571 9877 4580 9911
rect 4528 9868 4580 9877
rect 6644 9868 6696 9920
rect 6920 9868 6972 9920
rect 7196 9868 7248 9920
rect 7840 9868 7892 9920
rect 8024 9868 8076 9920
rect 9036 9868 9088 9920
rect 12532 9868 12584 9920
rect 12900 9868 12952 9920
rect 13912 9868 13964 9920
rect 16028 9868 16080 9920
rect 17224 9868 17276 9920
rect 19892 9868 19944 9920
rect 20720 9868 20772 9920
rect 21364 9936 21416 9988
rect 21548 9868 21600 9920
rect 23204 10072 23256 10124
rect 24400 10072 24452 10124
rect 24492 10072 24544 10124
rect 25596 10140 25648 10192
rect 26516 10140 26568 10192
rect 31668 10251 31720 10260
rect 31668 10217 31677 10251
rect 31677 10217 31711 10251
rect 31711 10217 31720 10251
rect 31668 10208 31720 10217
rect 32404 10208 32456 10260
rect 32680 10208 32732 10260
rect 32956 10251 33008 10260
rect 32956 10217 32965 10251
rect 32965 10217 32999 10251
rect 32999 10217 33008 10251
rect 32956 10208 33008 10217
rect 27160 10140 27212 10192
rect 27620 10140 27672 10192
rect 26792 10072 26844 10124
rect 29736 10140 29788 10192
rect 22652 10047 22704 10056
rect 22652 10013 22661 10047
rect 22661 10013 22695 10047
rect 22695 10013 22704 10047
rect 22652 10004 22704 10013
rect 23756 10004 23808 10056
rect 24768 9936 24820 9988
rect 25044 10004 25096 10056
rect 25688 9979 25740 9988
rect 25688 9945 25697 9979
rect 25697 9945 25731 9979
rect 25731 9945 25740 9979
rect 25688 9936 25740 9945
rect 26148 9979 26200 9988
rect 26148 9945 26157 9979
rect 26157 9945 26191 9979
rect 26191 9945 26200 9979
rect 26148 9936 26200 9945
rect 27620 10004 27672 10056
rect 28356 10004 28408 10056
rect 23756 9868 23808 9920
rect 25044 9868 25096 9920
rect 25872 9868 25924 9920
rect 26240 9911 26292 9920
rect 26240 9877 26249 9911
rect 26249 9877 26283 9911
rect 26283 9877 26292 9911
rect 26240 9868 26292 9877
rect 27160 9936 27212 9988
rect 27436 9979 27488 9988
rect 27436 9945 27445 9979
rect 27445 9945 27479 9979
rect 27479 9945 27488 9979
rect 27436 9936 27488 9945
rect 27528 9979 27580 9988
rect 27528 9945 27537 9979
rect 27537 9945 27571 9979
rect 27571 9945 27580 9979
rect 27528 9936 27580 9945
rect 28264 9936 28316 9988
rect 28908 10047 28960 10058
rect 28908 10013 28917 10047
rect 28917 10013 28951 10047
rect 28951 10013 28960 10047
rect 28908 10006 28960 10013
rect 30012 10004 30064 10056
rect 30748 10047 30800 10056
rect 30748 10013 30757 10047
rect 30757 10013 30791 10047
rect 30791 10013 30800 10047
rect 30748 10004 30800 10013
rect 27344 9868 27396 9920
rect 28080 9868 28132 9920
rect 31024 10115 31076 10124
rect 31024 10081 31033 10115
rect 31033 10081 31067 10115
rect 31067 10081 31076 10115
rect 31024 10072 31076 10081
rect 36544 10208 36596 10260
rect 32036 10072 32088 10124
rect 31944 10004 31996 10056
rect 32404 10047 32456 10056
rect 32404 10013 32413 10047
rect 32413 10013 32447 10047
rect 32447 10013 32456 10047
rect 32404 10004 32456 10013
rect 32772 10047 32824 10056
rect 32772 10013 32781 10047
rect 32781 10013 32815 10047
rect 32815 10013 32824 10047
rect 32772 10004 32824 10013
rect 33416 10047 33468 10056
rect 33416 10013 33425 10047
rect 33425 10013 33459 10047
rect 33459 10013 33468 10047
rect 33416 10004 33468 10013
rect 37004 10140 37056 10192
rect 34060 10072 34112 10124
rect 34612 10072 34664 10124
rect 33968 10004 34020 10056
rect 37464 10004 37516 10056
rect 39396 10004 39448 10056
rect 29736 9868 29788 9920
rect 29828 9911 29880 9920
rect 29828 9877 29837 9911
rect 29837 9877 29871 9911
rect 29871 9877 29880 9911
rect 29828 9868 29880 9877
rect 30012 9868 30064 9920
rect 30196 9868 30248 9920
rect 31392 9868 31444 9920
rect 31852 9868 31904 9920
rect 32864 9936 32916 9988
rect 35164 9979 35216 9988
rect 35164 9945 35173 9979
rect 35173 9945 35207 9979
rect 35207 9945 35216 9979
rect 35164 9936 35216 9945
rect 36452 9936 36504 9988
rect 33968 9911 34020 9920
rect 33968 9877 33977 9911
rect 33977 9877 34011 9911
rect 34011 9877 34020 9911
rect 33968 9868 34020 9877
rect 35348 9868 35400 9920
rect 37556 9868 37608 9920
rect 10472 9766 10524 9818
rect 10536 9766 10588 9818
rect 10600 9766 10652 9818
rect 10664 9766 10716 9818
rect 10728 9766 10780 9818
rect 19994 9766 20046 9818
rect 20058 9766 20110 9818
rect 20122 9766 20174 9818
rect 20186 9766 20238 9818
rect 20250 9766 20302 9818
rect 29516 9766 29568 9818
rect 29580 9766 29632 9818
rect 29644 9766 29696 9818
rect 29708 9766 29760 9818
rect 29772 9766 29824 9818
rect 39038 9766 39090 9818
rect 39102 9766 39154 9818
rect 39166 9766 39218 9818
rect 39230 9766 39282 9818
rect 39294 9766 39346 9818
rect 7104 9664 7156 9716
rect 13820 9664 13872 9716
rect 16120 9664 16172 9716
rect 16488 9664 16540 9716
rect 16856 9664 16908 9716
rect 1400 9528 1452 9580
rect 5540 9596 5592 9648
rect 6368 9596 6420 9648
rect 8760 9596 8812 9648
rect 9680 9596 9732 9648
rect 11152 9596 11204 9648
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 2412 9503 2464 9512
rect 2412 9469 2421 9503
rect 2421 9469 2455 9503
rect 2455 9469 2464 9503
rect 2412 9460 2464 9469
rect 4160 9460 4212 9512
rect 4252 9460 4304 9512
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 11980 9528 12032 9580
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 12716 9596 12768 9648
rect 13912 9528 13964 9580
rect 6276 9460 6328 9512
rect 6828 9460 6880 9512
rect 7380 9503 7432 9512
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 8116 9460 8168 9512
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9312 9460 9364 9469
rect 9588 9503 9640 9512
rect 9588 9469 9597 9503
rect 9597 9469 9631 9503
rect 9631 9469 9640 9503
rect 9588 9460 9640 9469
rect 9680 9460 9732 9512
rect 11612 9460 11664 9512
rect 11888 9460 11940 9512
rect 13176 9460 13228 9512
rect 14464 9528 14516 9580
rect 14648 9528 14700 9580
rect 8484 9392 8536 9444
rect 8760 9392 8812 9444
rect 10600 9392 10652 9444
rect 12072 9392 12124 9444
rect 12716 9392 12768 9444
rect 15108 9460 15160 9512
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 16212 9639 16264 9648
rect 16212 9605 16221 9639
rect 16221 9605 16255 9639
rect 16255 9605 16264 9639
rect 16212 9596 16264 9605
rect 17040 9596 17092 9648
rect 17776 9639 17828 9648
rect 17776 9605 17785 9639
rect 17785 9605 17819 9639
rect 17819 9605 17828 9639
rect 17776 9596 17828 9605
rect 17960 9664 18012 9716
rect 19892 9664 19944 9716
rect 20812 9664 20864 9716
rect 20352 9596 20404 9648
rect 16304 9528 16356 9580
rect 16488 9528 16540 9580
rect 16764 9528 16816 9580
rect 20444 9528 20496 9580
rect 20996 9528 21048 9580
rect 17592 9460 17644 9512
rect 17868 9460 17920 9512
rect 4528 9324 4580 9376
rect 5540 9324 5592 9376
rect 6092 9324 6144 9376
rect 7196 9324 7248 9376
rect 7564 9324 7616 9376
rect 8944 9324 8996 9376
rect 11704 9324 11756 9376
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 15476 9392 15528 9444
rect 16212 9392 16264 9444
rect 19708 9460 19760 9512
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 22652 9664 22704 9716
rect 26516 9664 26568 9716
rect 22560 9596 22612 9648
rect 21272 9528 21324 9537
rect 23940 9596 23992 9648
rect 24032 9639 24084 9648
rect 24032 9605 24041 9639
rect 24041 9605 24075 9639
rect 24075 9605 24084 9639
rect 24032 9596 24084 9605
rect 25320 9596 25372 9648
rect 23664 9528 23716 9580
rect 25136 9528 25188 9580
rect 25688 9528 25740 9580
rect 26792 9596 26844 9648
rect 27896 9639 27948 9648
rect 27896 9605 27905 9639
rect 27905 9605 27939 9639
rect 27939 9605 27948 9639
rect 27896 9596 27948 9605
rect 27988 9639 28040 9648
rect 27988 9605 27997 9639
rect 27997 9605 28031 9639
rect 28031 9605 28040 9639
rect 27988 9596 28040 9605
rect 22744 9503 22796 9512
rect 22744 9469 22753 9503
rect 22753 9469 22787 9503
rect 22787 9469 22796 9503
rect 22744 9460 22796 9469
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 18236 9324 18288 9376
rect 23756 9392 23808 9444
rect 26148 9392 26200 9444
rect 26700 9528 26752 9580
rect 27528 9460 27580 9512
rect 26516 9392 26568 9444
rect 27160 9392 27212 9444
rect 25320 9324 25372 9376
rect 25504 9367 25556 9376
rect 25504 9333 25513 9367
rect 25513 9333 25547 9367
rect 25547 9333 25556 9367
rect 25504 9324 25556 9333
rect 25596 9324 25648 9376
rect 26792 9324 26844 9376
rect 27436 9324 27488 9376
rect 27896 9460 27948 9512
rect 27712 9392 27764 9444
rect 29092 9664 29144 9716
rect 29460 9664 29512 9716
rect 29552 9664 29604 9716
rect 30288 9664 30340 9716
rect 29184 9596 29236 9648
rect 31024 9664 31076 9716
rect 31668 9664 31720 9716
rect 33048 9664 33100 9716
rect 28356 9460 28408 9512
rect 30012 9503 30064 9512
rect 30012 9469 30021 9503
rect 30021 9469 30055 9503
rect 30055 9469 30064 9503
rect 30012 9460 30064 9469
rect 31024 9460 31076 9512
rect 29184 9392 29236 9444
rect 33784 9596 33836 9648
rect 34520 9596 34572 9648
rect 31944 9528 31996 9580
rect 35624 9571 35676 9580
rect 35624 9537 35633 9571
rect 35633 9537 35667 9571
rect 35667 9537 35676 9571
rect 35624 9528 35676 9537
rect 32588 9503 32640 9512
rect 32588 9469 32597 9503
rect 32597 9469 32631 9503
rect 32631 9469 32640 9503
rect 32588 9460 32640 9469
rect 33232 9503 33284 9512
rect 33232 9469 33241 9503
rect 33241 9469 33275 9503
rect 33275 9469 33284 9503
rect 33232 9460 33284 9469
rect 36544 9596 36596 9648
rect 37464 9571 37516 9580
rect 37464 9537 37473 9571
rect 37473 9537 37507 9571
rect 37507 9537 37516 9571
rect 37464 9528 37516 9537
rect 38108 9571 38160 9580
rect 38108 9537 38117 9571
rect 38117 9537 38151 9571
rect 38151 9537 38160 9571
rect 38108 9528 38160 9537
rect 37924 9460 37976 9512
rect 31484 9324 31536 9376
rect 33324 9324 33376 9376
rect 38200 9367 38252 9376
rect 38200 9333 38209 9367
rect 38209 9333 38243 9367
rect 38243 9333 38252 9367
rect 38200 9324 38252 9333
rect 5711 9222 5763 9274
rect 5775 9222 5827 9274
rect 5839 9222 5891 9274
rect 5903 9222 5955 9274
rect 5967 9222 6019 9274
rect 15233 9222 15285 9274
rect 15297 9222 15349 9274
rect 15361 9222 15413 9274
rect 15425 9222 15477 9274
rect 15489 9222 15541 9274
rect 24755 9222 24807 9274
rect 24819 9222 24871 9274
rect 24883 9222 24935 9274
rect 24947 9222 24999 9274
rect 25011 9222 25063 9274
rect 34277 9222 34329 9274
rect 34341 9222 34393 9274
rect 34405 9222 34457 9274
rect 34469 9222 34521 9274
rect 34533 9222 34585 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 2964 9120 3016 9172
rect 4068 9120 4120 9172
rect 6000 9120 6052 9172
rect 7380 9120 7432 9172
rect 7748 9120 7800 9172
rect 8208 9120 8260 9172
rect 8392 9163 8444 9172
rect 8392 9129 8401 9163
rect 8401 9129 8435 9163
rect 8435 9129 8444 9163
rect 8392 9120 8444 9129
rect 9588 9120 9640 9172
rect 2412 9052 2464 9104
rect 2136 8984 2188 9036
rect 2596 8984 2648 9036
rect 3148 8984 3200 9036
rect 3700 8984 3752 9036
rect 6092 9052 6144 9104
rect 8944 9052 8996 9104
rect 14740 9120 14792 9172
rect 15568 9120 15620 9172
rect 4252 8984 4304 9036
rect 4804 8984 4856 9036
rect 7104 9027 7156 9036
rect 7104 8993 7113 9027
rect 7113 8993 7147 9027
rect 7147 8993 7156 9027
rect 7104 8984 7156 8993
rect 20 8916 72 8968
rect 3792 8916 3844 8968
rect 5632 8916 5684 8968
rect 7564 8916 7616 8968
rect 9680 8984 9732 9036
rect 10324 8984 10376 9036
rect 10968 8984 11020 9036
rect 11336 8984 11388 9036
rect 12532 9052 12584 9104
rect 7840 8959 7892 8968
rect 7840 8925 7850 8959
rect 7850 8925 7884 8959
rect 7884 8925 7892 8959
rect 7840 8916 7892 8925
rect 7932 8916 7984 8968
rect 8208 8959 8260 8968
rect 8208 8925 8222 8959
rect 8222 8925 8256 8959
rect 8256 8925 8260 8959
rect 8208 8916 8260 8925
rect 4988 8848 5040 8900
rect 6368 8848 6420 8900
rect 5080 8780 5132 8832
rect 6828 8780 6880 8832
rect 7196 8780 7248 8832
rect 7748 8780 7800 8832
rect 8024 8891 8076 8900
rect 8024 8857 8033 8891
rect 8033 8857 8067 8891
rect 8067 8857 8076 8891
rect 8024 8848 8076 8857
rect 9680 8848 9732 8900
rect 10416 8916 10468 8968
rect 10600 8848 10652 8900
rect 10784 8780 10836 8832
rect 11888 8848 11940 8900
rect 13452 9027 13504 9036
rect 13452 8993 13461 9027
rect 13461 8993 13495 9027
rect 13495 8993 13504 9027
rect 13452 8984 13504 8993
rect 14464 9052 14516 9104
rect 14832 9052 14884 9104
rect 13912 8984 13964 9036
rect 14188 8984 14240 9036
rect 14280 8916 14332 8968
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 12900 8848 12952 8900
rect 15108 8984 15160 9036
rect 14832 8959 14884 8968
rect 14832 8925 14835 8959
rect 14835 8925 14884 8959
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 15844 8984 15896 9036
rect 14832 8916 14884 8925
rect 13636 8780 13688 8832
rect 14740 8780 14792 8832
rect 15384 8848 15436 8900
rect 15752 8891 15804 8900
rect 15752 8857 15761 8891
rect 15761 8857 15795 8891
rect 15795 8857 15804 8891
rect 15752 8848 15804 8857
rect 15292 8780 15344 8832
rect 17592 8916 17644 8968
rect 18236 8916 18288 8968
rect 22376 9120 22428 9172
rect 25596 9120 25648 9172
rect 26240 9120 26292 9172
rect 26424 9120 26476 9172
rect 26608 9120 26660 9172
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 19340 8984 19392 9036
rect 20536 9027 20588 9036
rect 20536 8993 20545 9027
rect 20545 8993 20579 9027
rect 20579 8993 20588 9027
rect 20536 8984 20588 8993
rect 30748 9120 30800 9172
rect 31024 9120 31076 9172
rect 34704 9120 34756 9172
rect 35164 9120 35216 9172
rect 36176 9163 36228 9172
rect 36176 9129 36185 9163
rect 36185 9129 36219 9163
rect 36219 9129 36228 9163
rect 36176 9120 36228 9129
rect 38568 9163 38620 9172
rect 38568 9129 38577 9163
rect 38577 9129 38611 9163
rect 38611 9129 38620 9163
rect 38568 9120 38620 9129
rect 29276 9052 29328 9104
rect 30196 9052 30248 9104
rect 32588 9052 32640 9104
rect 34612 9052 34664 9104
rect 35624 9052 35676 9104
rect 23664 8984 23716 9036
rect 26424 8984 26476 9036
rect 26608 8984 26660 9036
rect 28540 8984 28592 9036
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 19984 8916 20036 8968
rect 21916 8916 21968 8968
rect 23480 8916 23532 8968
rect 26792 8916 26844 8968
rect 29552 8916 29604 8968
rect 17500 8891 17552 8900
rect 17500 8857 17509 8891
rect 17509 8857 17543 8891
rect 17543 8857 17552 8891
rect 17500 8848 17552 8857
rect 18604 8891 18656 8900
rect 18604 8857 18613 8891
rect 18613 8857 18647 8891
rect 18647 8857 18656 8891
rect 18604 8848 18656 8857
rect 18696 8780 18748 8832
rect 19432 8780 19484 8832
rect 20628 8780 20680 8832
rect 20812 8891 20864 8900
rect 20812 8857 20821 8891
rect 20821 8857 20855 8891
rect 20855 8857 20864 8891
rect 20812 8848 20864 8857
rect 24492 8848 24544 8900
rect 24860 8891 24912 8900
rect 24860 8857 24869 8891
rect 24869 8857 24903 8891
rect 24903 8857 24912 8891
rect 24860 8848 24912 8857
rect 29920 8984 29972 9036
rect 30012 8984 30064 9036
rect 31760 8984 31812 9036
rect 32772 8984 32824 9036
rect 30288 8916 30340 8968
rect 33600 8916 33652 8968
rect 33692 8959 33744 8968
rect 33692 8925 33701 8959
rect 33701 8925 33735 8959
rect 33735 8925 33744 8959
rect 33692 8916 33744 8925
rect 34888 8984 34940 9036
rect 35164 8984 35216 9036
rect 35348 9027 35400 9036
rect 35348 8993 35357 9027
rect 35357 8993 35391 9027
rect 35391 8993 35400 9027
rect 35348 8984 35400 8993
rect 35532 9027 35584 9036
rect 35532 8993 35541 9027
rect 35541 8993 35575 9027
rect 35575 8993 35584 9027
rect 35532 8984 35584 8993
rect 35900 8984 35952 9036
rect 35256 8959 35308 8968
rect 35256 8925 35265 8959
rect 35265 8925 35299 8959
rect 35299 8925 35308 8959
rect 35256 8916 35308 8925
rect 35624 8916 35676 8968
rect 29920 8891 29972 8900
rect 22468 8780 22520 8832
rect 26424 8780 26476 8832
rect 29920 8857 29929 8891
rect 29929 8857 29963 8891
rect 29963 8857 29972 8891
rect 29920 8848 29972 8857
rect 30196 8848 30248 8900
rect 30472 8848 30524 8900
rect 28908 8780 28960 8832
rect 30748 8780 30800 8832
rect 33784 8891 33836 8900
rect 33784 8857 33793 8891
rect 33793 8857 33827 8891
rect 33827 8857 33836 8891
rect 33784 8848 33836 8857
rect 34060 8823 34112 8832
rect 34060 8789 34069 8823
rect 34069 8789 34103 8823
rect 34103 8789 34112 8823
rect 34060 8780 34112 8789
rect 34888 8848 34940 8900
rect 36728 8848 36780 8900
rect 37096 8891 37148 8900
rect 37096 8857 37105 8891
rect 37105 8857 37139 8891
rect 37139 8857 37148 8891
rect 37096 8848 37148 8857
rect 37556 8848 37608 8900
rect 35624 8780 35676 8832
rect 10472 8678 10524 8730
rect 10536 8678 10588 8730
rect 10600 8678 10652 8730
rect 10664 8678 10716 8730
rect 10728 8678 10780 8730
rect 19994 8678 20046 8730
rect 20058 8678 20110 8730
rect 20122 8678 20174 8730
rect 20186 8678 20238 8730
rect 20250 8678 20302 8730
rect 29516 8678 29568 8730
rect 29580 8678 29632 8730
rect 29644 8678 29696 8730
rect 29708 8678 29760 8730
rect 29772 8678 29824 8730
rect 39038 8678 39090 8730
rect 39102 8678 39154 8730
rect 39166 8678 39218 8730
rect 39230 8678 39282 8730
rect 39294 8678 39346 8730
rect 3332 8576 3384 8628
rect 4252 8576 4304 8628
rect 6276 8576 6328 8628
rect 6828 8576 6880 8628
rect 8944 8576 8996 8628
rect 9496 8576 9548 8628
rect 4620 8508 4672 8560
rect 7472 8508 7524 8560
rect 8576 8551 8628 8560
rect 8576 8517 8585 8551
rect 8585 8517 8619 8551
rect 8619 8517 8628 8551
rect 8576 8508 8628 8517
rect 10140 8508 10192 8560
rect 11428 8576 11480 8628
rect 10784 8551 10836 8560
rect 10784 8517 10793 8551
rect 10793 8517 10827 8551
rect 10827 8517 10836 8551
rect 10784 8508 10836 8517
rect 940 8440 992 8492
rect 2780 8440 2832 8492
rect 3148 8440 3200 8492
rect 1952 8372 2004 8424
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 6828 8440 6880 8492
rect 7380 8440 7432 8492
rect 7932 8440 7984 8492
rect 11244 8440 11296 8492
rect 11428 8440 11480 8492
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 7196 8372 7248 8424
rect 8116 8372 8168 8424
rect 9772 8372 9824 8424
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12532 8576 12584 8628
rect 12072 8508 12124 8560
rect 13176 8551 13228 8560
rect 13176 8517 13185 8551
rect 13185 8517 13219 8551
rect 13219 8517 13228 8551
rect 13176 8508 13228 8517
rect 13912 8576 13964 8628
rect 14924 8576 14976 8628
rect 15384 8576 15436 8628
rect 15752 8576 15804 8628
rect 20812 8576 20864 8628
rect 22192 8576 22244 8628
rect 22468 8619 22520 8628
rect 22468 8585 22477 8619
rect 22477 8585 22511 8619
rect 22511 8585 22520 8619
rect 22468 8576 22520 8585
rect 23848 8576 23900 8628
rect 14280 8508 14332 8560
rect 17040 8508 17092 8560
rect 17132 8551 17184 8560
rect 17132 8517 17141 8551
rect 17141 8517 17175 8551
rect 17175 8517 17184 8551
rect 17132 8508 17184 8517
rect 17592 8508 17644 8560
rect 12624 8440 12676 8492
rect 14832 8440 14884 8492
rect 3332 8236 3384 8288
rect 5632 8236 5684 8288
rect 6828 8236 6880 8288
rect 9956 8236 10008 8288
rect 10784 8236 10836 8288
rect 13176 8372 13228 8424
rect 14556 8372 14608 8424
rect 15752 8440 15804 8492
rect 16672 8440 16724 8492
rect 16764 8440 16816 8492
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 14280 8304 14332 8356
rect 13268 8236 13320 8288
rect 15384 8372 15436 8424
rect 16396 8372 16448 8424
rect 24032 8508 24084 8560
rect 20352 8440 20404 8492
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 21548 8440 21600 8492
rect 15752 8304 15804 8356
rect 16028 8304 16080 8356
rect 18512 8304 18564 8356
rect 19432 8304 19484 8356
rect 19892 8372 19944 8424
rect 20536 8372 20588 8424
rect 20996 8372 21048 8424
rect 23020 8372 23072 8424
rect 24400 8440 24452 8492
rect 24860 8576 24912 8628
rect 25964 8576 26016 8628
rect 26240 8619 26292 8628
rect 26240 8585 26249 8619
rect 26249 8585 26283 8619
rect 26283 8585 26292 8619
rect 26240 8576 26292 8585
rect 24768 8508 24820 8560
rect 27436 8551 27488 8560
rect 27436 8517 27445 8551
rect 27445 8517 27479 8551
rect 27479 8517 27488 8551
rect 27436 8508 27488 8517
rect 28448 8508 28500 8560
rect 28908 8619 28960 8628
rect 28908 8585 28917 8619
rect 28917 8585 28951 8619
rect 28951 8585 28960 8619
rect 28908 8576 28960 8585
rect 29000 8576 29052 8628
rect 29828 8576 29880 8628
rect 29920 8576 29972 8628
rect 31852 8576 31904 8628
rect 32312 8619 32364 8628
rect 32312 8585 32321 8619
rect 32321 8585 32355 8619
rect 32355 8585 32364 8619
rect 32312 8576 32364 8585
rect 32496 8576 32548 8628
rect 32864 8576 32916 8628
rect 33416 8576 33468 8628
rect 34704 8576 34756 8628
rect 37924 8619 37976 8628
rect 37924 8585 37933 8619
rect 37933 8585 37967 8619
rect 37967 8585 37976 8619
rect 37924 8576 37976 8585
rect 30196 8508 30248 8560
rect 31024 8551 31076 8560
rect 31024 8517 31033 8551
rect 31033 8517 31067 8551
rect 31067 8517 31076 8551
rect 31024 8508 31076 8517
rect 31392 8508 31444 8560
rect 31668 8508 31720 8560
rect 33600 8508 33652 8560
rect 25780 8440 25832 8492
rect 28908 8440 28960 8492
rect 33324 8440 33376 8492
rect 25596 8372 25648 8424
rect 26516 8372 26568 8424
rect 26792 8372 26844 8424
rect 16672 8236 16724 8288
rect 17500 8236 17552 8288
rect 19616 8236 19668 8288
rect 19800 8236 19852 8288
rect 20260 8304 20312 8356
rect 25504 8304 25556 8356
rect 25688 8304 25740 8356
rect 25964 8304 26016 8356
rect 27896 8372 27948 8424
rect 30288 8372 30340 8424
rect 31208 8415 31260 8424
rect 31208 8381 31217 8415
rect 31217 8381 31251 8415
rect 31251 8381 31260 8415
rect 31208 8372 31260 8381
rect 32956 8415 33008 8424
rect 32956 8381 32965 8415
rect 32965 8381 32999 8415
rect 32999 8381 33008 8415
rect 32956 8372 33008 8381
rect 33876 8483 33928 8492
rect 33876 8449 33885 8483
rect 33885 8449 33919 8483
rect 33919 8449 33928 8483
rect 33876 8440 33928 8449
rect 34888 8483 34940 8492
rect 34888 8449 34897 8483
rect 34897 8449 34931 8483
rect 34931 8449 34940 8483
rect 34888 8440 34940 8449
rect 35440 8508 35492 8560
rect 28816 8304 28868 8356
rect 29000 8304 29052 8356
rect 29092 8304 29144 8356
rect 29552 8304 29604 8356
rect 34060 8415 34112 8424
rect 34060 8381 34069 8415
rect 34069 8381 34103 8415
rect 34103 8381 34112 8415
rect 34060 8372 34112 8381
rect 35164 8415 35216 8424
rect 35164 8381 35173 8415
rect 35173 8381 35207 8415
rect 35207 8381 35216 8415
rect 35164 8372 35216 8381
rect 35532 8372 35584 8424
rect 35992 8483 36044 8492
rect 35992 8449 36001 8483
rect 36001 8449 36035 8483
rect 36035 8449 36044 8483
rect 35992 8440 36044 8449
rect 37832 8483 37884 8492
rect 37832 8449 37841 8483
rect 37841 8449 37875 8483
rect 37875 8449 37884 8483
rect 37832 8440 37884 8449
rect 36912 8372 36964 8424
rect 33416 8304 33468 8356
rect 21456 8236 21508 8288
rect 25136 8236 25188 8288
rect 30196 8236 30248 8288
rect 31668 8236 31720 8288
rect 33048 8236 33100 8288
rect 33784 8236 33836 8288
rect 34060 8236 34112 8288
rect 34888 8236 34940 8288
rect 35164 8236 35216 8288
rect 35348 8304 35400 8356
rect 5711 8134 5763 8186
rect 5775 8134 5827 8186
rect 5839 8134 5891 8186
rect 5903 8134 5955 8186
rect 5967 8134 6019 8186
rect 15233 8134 15285 8186
rect 15297 8134 15349 8186
rect 15361 8134 15413 8186
rect 15425 8134 15477 8186
rect 15489 8134 15541 8186
rect 24755 8134 24807 8186
rect 24819 8134 24871 8186
rect 24883 8134 24935 8186
rect 24947 8134 24999 8186
rect 25011 8134 25063 8186
rect 34277 8134 34329 8186
rect 34341 8134 34393 8186
rect 34405 8134 34457 8186
rect 34469 8134 34521 8186
rect 34533 8134 34585 8186
rect 2964 8032 3016 8084
rect 3332 8032 3384 8084
rect 4436 8075 4488 8084
rect 4436 8041 4445 8075
rect 4445 8041 4479 8075
rect 4479 8041 4488 8075
rect 4436 8032 4488 8041
rect 3884 7964 3936 8016
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 4620 7896 4672 7948
rect 9036 8032 9088 8084
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 7104 7896 7156 7948
rect 7564 7896 7616 7948
rect 8852 7896 8904 7948
rect 10784 8032 10836 8084
rect 12348 7964 12400 8016
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 16304 8032 16356 8084
rect 17776 8032 17828 8084
rect 17960 8032 18012 8084
rect 18144 8032 18196 8084
rect 18972 8032 19024 8084
rect 14556 7964 14608 8016
rect 15844 7964 15896 8016
rect 10692 7896 10744 7948
rect 11060 7939 11112 7948
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 1952 7803 2004 7812
rect 1952 7769 1961 7803
rect 1961 7769 1995 7803
rect 1995 7769 2004 7803
rect 1952 7760 2004 7769
rect 2136 7803 2188 7812
rect 2136 7769 2177 7803
rect 2177 7769 2188 7803
rect 2136 7760 2188 7769
rect 2688 7760 2740 7812
rect 4344 7828 4396 7880
rect 5632 7828 5684 7880
rect 8576 7828 8628 7880
rect 9128 7828 9180 7880
rect 2412 7692 2464 7744
rect 4712 7760 4764 7812
rect 3884 7692 3936 7744
rect 7288 7760 7340 7812
rect 8484 7760 8536 7812
rect 13636 7828 13688 7880
rect 14556 7828 14608 7880
rect 15016 7828 15068 7880
rect 15200 7896 15252 7948
rect 15568 7896 15620 7948
rect 15752 7896 15804 7948
rect 19432 7964 19484 8016
rect 22284 8032 22336 8084
rect 23756 7964 23808 8016
rect 16764 7939 16816 7948
rect 16764 7905 16773 7939
rect 16773 7905 16807 7939
rect 16807 7905 16816 7939
rect 16764 7896 16816 7905
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 10968 7760 11020 7812
rect 11520 7760 11572 7812
rect 15752 7760 15804 7812
rect 16580 7760 16632 7812
rect 17500 7803 17552 7812
rect 17500 7769 17509 7803
rect 17509 7769 17543 7803
rect 17543 7769 17552 7803
rect 17500 7760 17552 7769
rect 17776 7828 17828 7880
rect 17960 7828 18012 7880
rect 23480 7896 23532 7948
rect 30196 8032 30248 8084
rect 23940 7964 23992 8016
rect 24768 7896 24820 7948
rect 24860 7896 24912 7948
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 19340 7828 19392 7880
rect 22192 7828 22244 7880
rect 23296 7828 23348 7880
rect 24952 7828 25004 7880
rect 18604 7803 18656 7812
rect 18604 7769 18613 7803
rect 18613 7769 18647 7803
rect 18647 7769 18656 7803
rect 18604 7760 18656 7769
rect 18788 7760 18840 7812
rect 20720 7760 20772 7812
rect 5080 7692 5132 7744
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 9588 7735 9640 7744
rect 9588 7701 9597 7735
rect 9597 7701 9631 7735
rect 9631 7701 9640 7735
rect 9588 7692 9640 7701
rect 13176 7692 13228 7744
rect 14280 7692 14332 7744
rect 14464 7692 14516 7744
rect 17960 7692 18012 7744
rect 19616 7692 19668 7744
rect 20260 7692 20312 7744
rect 20444 7692 20496 7744
rect 23940 7760 23992 7812
rect 24676 7760 24728 7812
rect 25136 7760 25188 7812
rect 25228 7760 25280 7812
rect 25504 7760 25556 7812
rect 21548 7735 21600 7744
rect 21548 7701 21557 7735
rect 21557 7701 21591 7735
rect 21591 7701 21600 7735
rect 21548 7692 21600 7701
rect 22652 7692 22704 7744
rect 23848 7692 23900 7744
rect 25320 7692 25372 7744
rect 25596 7692 25648 7744
rect 26056 7896 26108 7948
rect 26424 7896 26476 7948
rect 29092 7964 29144 8016
rect 31392 7964 31444 8016
rect 33324 8032 33376 8084
rect 34060 8032 34112 8084
rect 34520 8032 34572 8084
rect 34152 7964 34204 8016
rect 35808 7964 35860 8016
rect 37740 8007 37792 8016
rect 37740 7973 37749 8007
rect 37749 7973 37783 8007
rect 37783 7973 37792 8007
rect 37740 7964 37792 7973
rect 25872 7828 25924 7880
rect 26608 7828 26660 7880
rect 26792 7871 26844 7880
rect 26792 7837 26801 7871
rect 26801 7837 26835 7871
rect 26835 7837 26844 7871
rect 26792 7828 26844 7837
rect 28816 7871 28868 7880
rect 28816 7837 28825 7871
rect 28825 7837 28859 7871
rect 28859 7837 28868 7871
rect 28816 7828 28868 7837
rect 29000 7896 29052 7948
rect 30012 7896 30064 7948
rect 31760 7896 31812 7948
rect 33232 7896 33284 7948
rect 33968 7896 34020 7948
rect 25964 7803 26016 7812
rect 25964 7769 25973 7803
rect 25973 7769 26007 7803
rect 26007 7769 26016 7803
rect 25964 7760 26016 7769
rect 26056 7803 26108 7812
rect 26056 7769 26065 7803
rect 26065 7769 26099 7803
rect 26099 7769 26108 7803
rect 26056 7760 26108 7769
rect 26332 7735 26384 7744
rect 26332 7701 26341 7735
rect 26341 7701 26375 7735
rect 26375 7701 26384 7735
rect 26332 7692 26384 7701
rect 28724 7692 28776 7744
rect 28908 7692 28960 7744
rect 29092 7692 29144 7744
rect 31300 7692 31352 7744
rect 31668 7760 31720 7812
rect 32956 7760 33008 7812
rect 34704 7828 34756 7880
rect 35164 7939 35216 7948
rect 35164 7905 35173 7939
rect 35173 7905 35207 7939
rect 35207 7905 35216 7939
rect 35164 7896 35216 7905
rect 35900 7896 35952 7948
rect 35348 7871 35400 7880
rect 35348 7837 35357 7871
rect 35357 7837 35391 7871
rect 35391 7837 35400 7871
rect 35348 7828 35400 7837
rect 37004 7896 37056 7948
rect 37372 7828 37424 7880
rect 36176 7760 36228 7812
rect 36268 7803 36320 7812
rect 36268 7769 36277 7803
rect 36277 7769 36311 7803
rect 36311 7769 36320 7803
rect 36268 7760 36320 7769
rect 38660 7803 38712 7812
rect 38660 7769 38669 7803
rect 38669 7769 38703 7803
rect 38703 7769 38712 7803
rect 38660 7760 38712 7769
rect 35532 7735 35584 7744
rect 35532 7701 35541 7735
rect 35541 7701 35575 7735
rect 35575 7701 35584 7735
rect 35532 7692 35584 7701
rect 10472 7590 10524 7642
rect 10536 7590 10588 7642
rect 10600 7590 10652 7642
rect 10664 7590 10716 7642
rect 10728 7590 10780 7642
rect 19994 7590 20046 7642
rect 20058 7590 20110 7642
rect 20122 7590 20174 7642
rect 20186 7590 20238 7642
rect 20250 7590 20302 7642
rect 29516 7590 29568 7642
rect 29580 7590 29632 7642
rect 29644 7590 29696 7642
rect 29708 7590 29760 7642
rect 29772 7590 29824 7642
rect 39038 7590 39090 7642
rect 39102 7590 39154 7642
rect 39166 7590 39218 7642
rect 39230 7590 39282 7642
rect 39294 7590 39346 7642
rect 3332 7531 3384 7540
rect 3332 7497 3341 7531
rect 3341 7497 3375 7531
rect 3375 7497 3384 7531
rect 3332 7488 3384 7497
rect 4436 7488 4488 7540
rect 4804 7488 4856 7540
rect 7564 7488 7616 7540
rect 7656 7488 7708 7540
rect 2412 7420 2464 7472
rect 3608 7420 3660 7472
rect 1676 7352 1728 7404
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 3056 7395 3108 7404
rect 3056 7361 3065 7395
rect 3065 7361 3099 7395
rect 3099 7361 3108 7395
rect 3056 7352 3108 7361
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 6460 7420 6512 7472
rect 3148 7352 3200 7361
rect 3608 7284 3660 7336
rect 4436 7352 4488 7404
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 7380 7420 7432 7472
rect 15016 7488 15068 7540
rect 17040 7488 17092 7540
rect 18328 7488 18380 7540
rect 10416 7420 10468 7472
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 10876 7352 10928 7404
rect 11796 7352 11848 7404
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 5816 7327 5868 7336
rect 5816 7293 5825 7327
rect 5825 7293 5859 7327
rect 5859 7293 5868 7327
rect 5816 7284 5868 7293
rect 9128 7284 9180 7336
rect 9312 7284 9364 7336
rect 11244 7284 11296 7336
rect 12716 7420 12768 7472
rect 12992 7420 13044 7472
rect 14464 7420 14516 7472
rect 14740 7420 14792 7472
rect 16764 7420 16816 7472
rect 16948 7420 17000 7472
rect 21548 7488 21600 7540
rect 23388 7531 23440 7540
rect 23388 7497 23397 7531
rect 23397 7497 23431 7531
rect 23431 7497 23440 7531
rect 23388 7488 23440 7497
rect 24124 7488 24176 7540
rect 25688 7488 25740 7540
rect 25872 7488 25924 7540
rect 26976 7488 27028 7540
rect 27344 7488 27396 7540
rect 28172 7488 28224 7540
rect 12808 7352 12860 7404
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 2780 7216 2832 7268
rect 5080 7148 5132 7200
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 5632 7148 5684 7200
rect 6276 7148 6328 7200
rect 6552 7148 6604 7200
rect 6828 7148 6880 7200
rect 12072 7216 12124 7268
rect 12256 7216 12308 7268
rect 12532 7284 12584 7336
rect 13728 7352 13780 7404
rect 17316 7352 17368 7404
rect 18604 7352 18656 7404
rect 13452 7284 13504 7336
rect 17960 7284 18012 7336
rect 18880 7420 18932 7472
rect 20996 7420 21048 7472
rect 22468 7420 22520 7472
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 9588 7148 9640 7200
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 13820 7148 13872 7200
rect 14280 7148 14332 7200
rect 18144 7216 18196 7268
rect 20812 7284 20864 7336
rect 21456 7284 21508 7336
rect 22744 7395 22796 7404
rect 22744 7361 22753 7395
rect 22753 7361 22787 7395
rect 22787 7361 22796 7395
rect 22744 7352 22796 7361
rect 23296 7420 23348 7472
rect 23756 7395 23808 7404
rect 23756 7361 23765 7395
rect 23765 7361 23799 7395
rect 23799 7361 23808 7395
rect 23756 7352 23808 7361
rect 24492 7352 24544 7404
rect 25228 7420 25280 7472
rect 25504 7463 25556 7472
rect 25504 7429 25513 7463
rect 25513 7429 25547 7463
rect 25547 7429 25556 7463
rect 25504 7420 25556 7429
rect 27988 7420 28040 7472
rect 24860 7284 24912 7336
rect 25964 7352 26016 7404
rect 28356 7352 28408 7404
rect 29000 7420 29052 7472
rect 29368 7420 29420 7472
rect 31024 7488 31076 7540
rect 32404 7488 32456 7540
rect 32680 7488 32732 7540
rect 35256 7488 35308 7540
rect 34060 7463 34112 7472
rect 34060 7429 34069 7463
rect 34069 7429 34103 7463
rect 34103 7429 34112 7463
rect 34060 7420 34112 7429
rect 36176 7488 36228 7540
rect 36912 7531 36964 7540
rect 36912 7497 36921 7531
rect 36921 7497 36955 7531
rect 36955 7497 36964 7531
rect 36912 7488 36964 7497
rect 37188 7488 37240 7540
rect 31760 7352 31812 7404
rect 32680 7395 32732 7404
rect 32680 7361 32689 7395
rect 32689 7361 32723 7395
rect 32723 7361 32732 7395
rect 32680 7352 32732 7361
rect 33232 7352 33284 7404
rect 35992 7420 36044 7472
rect 25136 7284 25188 7336
rect 26792 7284 26844 7336
rect 16396 7148 16448 7200
rect 17132 7148 17184 7200
rect 17408 7148 17460 7200
rect 17868 7148 17920 7200
rect 21088 7148 21140 7200
rect 21180 7148 21232 7200
rect 24860 7191 24912 7200
rect 24860 7157 24869 7191
rect 24869 7157 24903 7191
rect 24903 7157 24912 7191
rect 24860 7148 24912 7157
rect 25780 7216 25832 7268
rect 27804 7284 27856 7336
rect 30288 7284 30340 7336
rect 31208 7284 31260 7336
rect 31576 7327 31628 7336
rect 31576 7293 31585 7327
rect 31585 7293 31619 7327
rect 31619 7293 31628 7327
rect 31576 7284 31628 7293
rect 32404 7284 32456 7336
rect 34704 7284 34756 7336
rect 25964 7148 26016 7200
rect 31392 7216 31444 7268
rect 37740 7284 37792 7336
rect 30288 7148 30340 7200
rect 31668 7148 31720 7200
rect 36728 7148 36780 7200
rect 5711 7046 5763 7098
rect 5775 7046 5827 7098
rect 5839 7046 5891 7098
rect 5903 7046 5955 7098
rect 5967 7046 6019 7098
rect 15233 7046 15285 7098
rect 15297 7046 15349 7098
rect 15361 7046 15413 7098
rect 15425 7046 15477 7098
rect 15489 7046 15541 7098
rect 24755 7046 24807 7098
rect 24819 7046 24871 7098
rect 24883 7046 24935 7098
rect 24947 7046 24999 7098
rect 25011 7046 25063 7098
rect 34277 7046 34329 7098
rect 34341 7046 34393 7098
rect 34405 7046 34457 7098
rect 34469 7046 34521 7098
rect 34533 7046 34585 7098
rect 2964 6944 3016 6996
rect 11704 6944 11756 6996
rect 12072 6944 12124 6996
rect 14740 6944 14792 6996
rect 15108 6944 15160 6996
rect 4436 6876 4488 6928
rect 1860 6808 1912 6860
rect 4344 6808 4396 6860
rect 12900 6876 12952 6928
rect 13636 6876 13688 6928
rect 14280 6876 14332 6928
rect 15384 6876 15436 6928
rect 15752 6876 15804 6928
rect 15936 6944 15988 6996
rect 17132 6944 17184 6996
rect 16672 6876 16724 6928
rect 18328 6944 18380 6996
rect 20812 6944 20864 6996
rect 21088 6987 21140 6996
rect 21088 6953 21097 6987
rect 21097 6953 21131 6987
rect 21131 6953 21140 6987
rect 21088 6944 21140 6953
rect 25228 6944 25280 6996
rect 26148 6944 26200 6996
rect 26976 6944 27028 6996
rect 27160 6944 27212 6996
rect 29000 6944 29052 6996
rect 31668 6944 31720 6996
rect 35992 6944 36044 6996
rect 36084 6944 36136 6996
rect 4804 6808 4856 6860
rect 6460 6808 6512 6860
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 10968 6808 11020 6860
rect 13728 6808 13780 6860
rect 16396 6808 16448 6860
rect 18236 6808 18288 6860
rect 18696 6808 18748 6860
rect 19340 6876 19392 6928
rect 20444 6851 20496 6860
rect 20444 6817 20453 6851
rect 20453 6817 20487 6851
rect 20487 6817 20496 6851
rect 20444 6808 20496 6817
rect 26608 6876 26660 6928
rect 23664 6808 23716 6860
rect 25136 6851 25188 6860
rect 25136 6817 25145 6851
rect 25145 6817 25179 6851
rect 25179 6817 25188 6851
rect 25136 6808 25188 6817
rect 25412 6808 25464 6860
rect 4436 6740 4488 6792
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 9772 6740 9824 6792
rect 10140 6740 10192 6792
rect 12440 6740 12492 6792
rect 12992 6740 13044 6792
rect 14004 6740 14056 6792
rect 15016 6740 15068 6792
rect 19524 6740 19576 6792
rect 20536 6740 20588 6792
rect 21088 6783 21140 6792
rect 21088 6749 21097 6783
rect 21097 6749 21131 6783
rect 21131 6749 21140 6783
rect 21088 6740 21140 6749
rect 1952 6672 2004 6724
rect 2136 6672 2188 6724
rect 2412 6672 2464 6724
rect 2596 6672 2648 6724
rect 2872 6672 2924 6724
rect 4160 6672 4212 6724
rect 4252 6672 4304 6724
rect 2320 6604 2372 6656
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 4068 6604 4120 6656
rect 6460 6672 6512 6724
rect 5540 6604 5592 6656
rect 7012 6672 7064 6724
rect 8392 6715 8444 6724
rect 8392 6681 8401 6715
rect 8401 6681 8435 6715
rect 8435 6681 8444 6715
rect 8392 6672 8444 6681
rect 11244 6672 11296 6724
rect 11336 6715 11388 6724
rect 11336 6681 11345 6715
rect 11345 6681 11379 6715
rect 11379 6681 11388 6715
rect 11336 6672 11388 6681
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 9864 6647 9916 6656
rect 9864 6613 9873 6647
rect 9873 6613 9907 6647
rect 9907 6613 9916 6647
rect 9864 6604 9916 6613
rect 15384 6672 15436 6724
rect 15476 6672 15528 6724
rect 16948 6672 17000 6724
rect 17500 6672 17552 6724
rect 18788 6715 18840 6724
rect 18788 6681 18797 6715
rect 18797 6681 18831 6715
rect 18831 6681 18840 6715
rect 18788 6672 18840 6681
rect 19708 6672 19760 6724
rect 20628 6672 20680 6724
rect 27528 6740 27580 6792
rect 27620 6783 27672 6792
rect 27620 6749 27629 6783
rect 27629 6749 27663 6783
rect 27663 6749 27672 6783
rect 27620 6740 27672 6749
rect 27804 6783 27856 6792
rect 27804 6749 27811 6783
rect 27811 6749 27856 6783
rect 27804 6740 27856 6749
rect 27988 6783 28040 6792
rect 27988 6749 27997 6783
rect 27997 6749 28031 6783
rect 28031 6749 28040 6783
rect 27988 6740 28040 6749
rect 28264 6876 28316 6928
rect 31392 6876 31444 6928
rect 31484 6876 31536 6928
rect 34888 6876 34940 6928
rect 30288 6808 30340 6860
rect 30748 6808 30800 6860
rect 28264 6740 28316 6792
rect 29276 6740 29328 6792
rect 31300 6808 31352 6860
rect 22928 6672 22980 6724
rect 15936 6604 15988 6656
rect 21456 6647 21508 6656
rect 21456 6613 21465 6647
rect 21465 6613 21499 6647
rect 21499 6613 21508 6647
rect 21456 6604 21508 6613
rect 25412 6715 25464 6724
rect 25412 6681 25421 6715
rect 25421 6681 25455 6715
rect 25455 6681 25464 6715
rect 25412 6672 25464 6681
rect 27344 6672 27396 6724
rect 28172 6604 28224 6656
rect 28264 6647 28316 6656
rect 28264 6613 28273 6647
rect 28273 6613 28307 6647
rect 28307 6613 28316 6647
rect 28264 6604 28316 6613
rect 30932 6672 30984 6724
rect 29920 6647 29972 6656
rect 29920 6613 29929 6647
rect 29929 6613 29963 6647
rect 29963 6613 29972 6647
rect 29920 6604 29972 6613
rect 30472 6647 30524 6656
rect 30472 6613 30481 6647
rect 30481 6613 30515 6647
rect 30515 6613 30524 6647
rect 30472 6604 30524 6613
rect 31484 6740 31536 6792
rect 31668 6783 31720 6792
rect 31668 6749 31677 6783
rect 31677 6749 31711 6783
rect 31711 6749 31720 6783
rect 31668 6740 31720 6749
rect 31852 6783 31904 6792
rect 31852 6749 31861 6783
rect 31861 6749 31895 6783
rect 31895 6749 31904 6783
rect 31852 6740 31904 6749
rect 32036 6783 32088 6792
rect 32036 6749 32045 6783
rect 32045 6749 32079 6783
rect 32079 6749 32088 6783
rect 32036 6740 32088 6749
rect 32680 6783 32732 6792
rect 32680 6749 32689 6783
rect 32689 6749 32723 6783
rect 32723 6749 32732 6783
rect 32680 6740 32732 6749
rect 37740 6808 37792 6860
rect 32772 6672 32824 6724
rect 33508 6715 33560 6724
rect 33508 6681 33517 6715
rect 33517 6681 33551 6715
rect 33551 6681 33560 6715
rect 33508 6672 33560 6681
rect 34060 6783 34112 6792
rect 34060 6749 34069 6783
rect 34069 6749 34103 6783
rect 34103 6749 34112 6783
rect 34060 6740 34112 6749
rect 34704 6740 34756 6792
rect 35808 6740 35860 6792
rect 35992 6740 36044 6792
rect 36084 6783 36136 6792
rect 36084 6749 36093 6783
rect 36093 6749 36127 6783
rect 36127 6749 36136 6783
rect 36084 6740 36136 6749
rect 36820 6783 36872 6792
rect 36820 6749 36829 6783
rect 36829 6749 36863 6783
rect 36863 6749 36872 6783
rect 36820 6740 36872 6749
rect 37372 6672 37424 6724
rect 34888 6647 34940 6656
rect 34888 6613 34897 6647
rect 34897 6613 34931 6647
rect 34931 6613 34940 6647
rect 34888 6604 34940 6613
rect 35256 6647 35308 6656
rect 35256 6613 35265 6647
rect 35265 6613 35299 6647
rect 35299 6613 35308 6647
rect 35256 6604 35308 6613
rect 37832 6604 37884 6656
rect 38568 6647 38620 6656
rect 38568 6613 38577 6647
rect 38577 6613 38611 6647
rect 38611 6613 38620 6647
rect 38568 6604 38620 6613
rect 10472 6502 10524 6554
rect 10536 6502 10588 6554
rect 10600 6502 10652 6554
rect 10664 6502 10716 6554
rect 10728 6502 10780 6554
rect 19994 6502 20046 6554
rect 20058 6502 20110 6554
rect 20122 6502 20174 6554
rect 20186 6502 20238 6554
rect 20250 6502 20302 6554
rect 29516 6502 29568 6554
rect 29580 6502 29632 6554
rect 29644 6502 29696 6554
rect 29708 6502 29760 6554
rect 29772 6502 29824 6554
rect 39038 6502 39090 6554
rect 39102 6502 39154 6554
rect 39166 6502 39218 6554
rect 39230 6502 39282 6554
rect 39294 6502 39346 6554
rect 3424 6400 3476 6452
rect 4252 6400 4304 6452
rect 3332 6332 3384 6384
rect 3976 6375 4028 6384
rect 3976 6341 3985 6375
rect 3985 6341 4019 6375
rect 4019 6341 4028 6375
rect 3976 6332 4028 6341
rect 4436 6332 4488 6384
rect 6460 6332 6512 6384
rect 6920 6400 6972 6452
rect 8024 6400 8076 6452
rect 10232 6400 10284 6452
rect 10784 6400 10836 6452
rect 12532 6443 12584 6452
rect 12532 6409 12541 6443
rect 12541 6409 12575 6443
rect 12575 6409 12584 6443
rect 12532 6400 12584 6409
rect 8300 6332 8352 6384
rect 13544 6400 13596 6452
rect 17224 6400 17276 6452
rect 17960 6400 18012 6452
rect 22560 6400 22612 6452
rect 22836 6400 22888 6452
rect 13360 6332 13412 6384
rect 940 6264 992 6316
rect 6368 6264 6420 6316
rect 2688 6196 2740 6248
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 3700 6239 3752 6248
rect 1584 6128 1636 6180
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 3700 6196 3752 6205
rect 3424 6128 3476 6180
rect 4068 6196 4120 6248
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7104 6264 7156 6316
rect 9128 6264 9180 6316
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 11244 6264 11296 6316
rect 12716 6264 12768 6316
rect 13820 6332 13872 6384
rect 15108 6332 15160 6384
rect 15844 6332 15896 6384
rect 18512 6375 18564 6384
rect 18512 6341 18521 6375
rect 18521 6341 18555 6375
rect 18555 6341 18564 6375
rect 18512 6332 18564 6341
rect 19800 6332 19852 6384
rect 20260 6332 20312 6384
rect 20628 6332 20680 6384
rect 20812 6375 20864 6384
rect 20812 6341 20821 6375
rect 20821 6341 20855 6375
rect 20855 6341 20864 6375
rect 20812 6332 20864 6341
rect 17500 6264 17552 6316
rect 23296 6332 23348 6384
rect 24216 6332 24268 6384
rect 24768 6332 24820 6384
rect 25504 6375 25556 6384
rect 25504 6341 25513 6375
rect 25513 6341 25547 6375
rect 25547 6341 25556 6375
rect 25504 6332 25556 6341
rect 27528 6400 27580 6452
rect 30288 6400 30340 6452
rect 31760 6400 31812 6452
rect 27896 6332 27948 6384
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 7012 6196 7064 6248
rect 1860 6060 1912 6112
rect 4528 6060 4580 6112
rect 7564 6128 7616 6180
rect 9312 6128 9364 6180
rect 12072 6128 12124 6180
rect 13084 6196 13136 6248
rect 13912 6239 13964 6248
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 14464 6196 14516 6248
rect 14556 6128 14608 6180
rect 5448 6060 5500 6112
rect 10508 6060 10560 6112
rect 10784 6060 10836 6112
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 13636 6060 13688 6112
rect 17868 6196 17920 6248
rect 16028 6128 16080 6180
rect 18972 6196 19024 6248
rect 19708 6196 19760 6248
rect 20352 6196 20404 6248
rect 20812 6196 20864 6248
rect 16580 6060 16632 6112
rect 20536 6128 20588 6180
rect 22284 6196 22336 6248
rect 22744 6264 22796 6316
rect 22100 6128 22152 6180
rect 23572 6196 23624 6248
rect 23020 6128 23072 6180
rect 25780 6264 25832 6316
rect 26148 6264 26200 6316
rect 25136 6196 25188 6248
rect 29920 6332 29972 6384
rect 31392 6332 31444 6384
rect 32680 6375 32732 6384
rect 32680 6341 32689 6375
rect 32689 6341 32723 6375
rect 32723 6341 32732 6375
rect 32680 6332 32732 6341
rect 31300 6264 31352 6316
rect 32496 6264 32548 6316
rect 26516 6128 26568 6180
rect 29368 6196 29420 6248
rect 32680 6196 32732 6248
rect 33048 6196 33100 6248
rect 33876 6375 33928 6384
rect 33876 6341 33885 6375
rect 33885 6341 33919 6375
rect 33919 6341 33928 6375
rect 33876 6332 33928 6341
rect 34152 6443 34204 6452
rect 34152 6409 34161 6443
rect 34161 6409 34195 6443
rect 34195 6409 34204 6443
rect 34152 6400 34204 6409
rect 37096 6400 37148 6452
rect 38476 6400 38528 6452
rect 36544 6332 36596 6384
rect 33968 6307 34020 6316
rect 33968 6273 33977 6307
rect 33977 6273 34011 6307
rect 34011 6273 34020 6307
rect 33968 6264 34020 6273
rect 36176 6264 36228 6316
rect 34244 6196 34296 6248
rect 19892 6060 19944 6112
rect 22192 6060 22244 6112
rect 24768 6060 24820 6112
rect 26240 6060 26292 6112
rect 29092 6060 29144 6112
rect 30104 6060 30156 6112
rect 31300 6060 31352 6112
rect 32680 6060 32732 6112
rect 32772 6060 32824 6112
rect 34152 6060 34204 6112
rect 34888 6239 34940 6248
rect 34888 6205 34897 6239
rect 34897 6205 34931 6239
rect 34931 6205 34940 6239
rect 34888 6196 34940 6205
rect 35624 6196 35676 6248
rect 37924 6196 37976 6248
rect 35992 6128 36044 6180
rect 35900 6060 35952 6112
rect 5711 5958 5763 6010
rect 5775 5958 5827 6010
rect 5839 5958 5891 6010
rect 5903 5958 5955 6010
rect 5967 5958 6019 6010
rect 15233 5958 15285 6010
rect 15297 5958 15349 6010
rect 15361 5958 15413 6010
rect 15425 5958 15477 6010
rect 15489 5958 15541 6010
rect 24755 5958 24807 6010
rect 24819 5958 24871 6010
rect 24883 5958 24935 6010
rect 24947 5958 24999 6010
rect 25011 5958 25063 6010
rect 34277 5958 34329 6010
rect 34341 5958 34393 6010
rect 34405 5958 34457 6010
rect 34469 5958 34521 6010
rect 34533 5958 34585 6010
rect 1952 5856 2004 5908
rect 2320 5720 2372 5772
rect 1584 5652 1636 5704
rect 3240 5584 3292 5636
rect 5264 5856 5316 5908
rect 7564 5856 7616 5908
rect 8300 5856 8352 5908
rect 8852 5856 8904 5908
rect 6276 5788 6328 5840
rect 6828 5788 6880 5840
rect 8116 5788 8168 5840
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 12992 5856 13044 5908
rect 13728 5856 13780 5908
rect 14464 5899 14516 5908
rect 14464 5865 14473 5899
rect 14473 5865 14507 5899
rect 14507 5865 14516 5899
rect 14464 5856 14516 5865
rect 14556 5856 14608 5908
rect 15752 5856 15804 5908
rect 17776 5856 17828 5908
rect 19616 5856 19668 5908
rect 20628 5856 20680 5908
rect 11980 5788 12032 5840
rect 14832 5788 14884 5840
rect 3700 5720 3752 5772
rect 4528 5652 4580 5704
rect 6552 5652 6604 5704
rect 8392 5720 8444 5772
rect 11060 5720 11112 5772
rect 11336 5652 11388 5704
rect 3976 5516 4028 5568
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 4896 5627 4948 5636
rect 4896 5593 4905 5627
rect 4905 5593 4939 5627
rect 4939 5593 4948 5627
rect 4896 5584 4948 5593
rect 6184 5584 6236 5636
rect 6644 5584 6696 5636
rect 11796 5584 11848 5636
rect 13544 5584 13596 5636
rect 14924 5763 14976 5772
rect 14924 5729 14933 5763
rect 14933 5729 14967 5763
rect 14967 5729 14976 5763
rect 14924 5720 14976 5729
rect 18144 5831 18196 5840
rect 18144 5797 18153 5831
rect 18153 5797 18187 5831
rect 18187 5797 18196 5831
rect 18144 5788 18196 5797
rect 15936 5763 15988 5772
rect 15936 5729 15945 5763
rect 15945 5729 15979 5763
rect 15979 5729 15988 5763
rect 15936 5720 15988 5729
rect 19708 5788 19760 5840
rect 20812 5788 20864 5840
rect 18696 5763 18748 5772
rect 18696 5729 18705 5763
rect 18705 5729 18739 5763
rect 18739 5729 18748 5763
rect 18696 5720 18748 5729
rect 19892 5720 19944 5772
rect 23020 5856 23072 5908
rect 23204 5899 23256 5908
rect 23204 5865 23213 5899
rect 23213 5865 23247 5899
rect 23247 5865 23256 5899
rect 23204 5856 23256 5865
rect 24584 5856 24636 5908
rect 25412 5856 25464 5908
rect 26332 5856 26384 5908
rect 26056 5788 26108 5840
rect 26424 5788 26476 5840
rect 30012 5788 30064 5840
rect 30104 5788 30156 5840
rect 25136 5720 25188 5772
rect 25596 5763 25648 5772
rect 14096 5652 14148 5704
rect 14556 5652 14608 5704
rect 15476 5652 15528 5704
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 17316 5652 17368 5704
rect 18328 5652 18380 5704
rect 19340 5652 19392 5704
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 20628 5695 20680 5704
rect 20628 5661 20637 5695
rect 20637 5661 20671 5695
rect 20671 5661 20680 5695
rect 20628 5652 20680 5661
rect 21088 5652 21140 5704
rect 5172 5516 5224 5568
rect 9772 5516 9824 5568
rect 11428 5516 11480 5568
rect 12072 5516 12124 5568
rect 13636 5516 13688 5568
rect 14740 5516 14792 5568
rect 16028 5584 16080 5636
rect 15476 5516 15528 5568
rect 17316 5516 17368 5568
rect 17960 5516 18012 5568
rect 19064 5516 19116 5568
rect 21180 5584 21232 5636
rect 21640 5584 21692 5636
rect 22376 5584 22428 5636
rect 22560 5516 22612 5568
rect 25596 5729 25605 5763
rect 25605 5729 25639 5763
rect 25639 5729 25648 5763
rect 25596 5720 25648 5729
rect 25964 5720 26016 5772
rect 26884 5720 26936 5772
rect 27068 5763 27120 5772
rect 27068 5729 27077 5763
rect 27077 5729 27111 5763
rect 27111 5729 27120 5763
rect 27068 5720 27120 5729
rect 27804 5720 27856 5772
rect 25320 5652 25372 5704
rect 26792 5695 26844 5704
rect 26792 5661 26801 5695
rect 26801 5661 26835 5695
rect 26835 5661 26844 5695
rect 26792 5652 26844 5661
rect 27436 5652 27488 5704
rect 27620 5652 27672 5704
rect 27988 5652 28040 5704
rect 28080 5695 28132 5704
rect 28080 5661 28089 5695
rect 28089 5661 28123 5695
rect 28123 5661 28132 5695
rect 28080 5652 28132 5661
rect 24768 5584 24820 5636
rect 26700 5584 26752 5636
rect 27528 5584 27580 5636
rect 28540 5720 28592 5772
rect 29920 5720 29972 5772
rect 30748 5788 30800 5840
rect 34888 5856 34940 5908
rect 35348 5856 35400 5908
rect 32404 5788 32456 5840
rect 30380 5720 30432 5772
rect 30932 5720 30984 5772
rect 32036 5720 32088 5772
rect 33508 5720 33560 5772
rect 28448 5652 28500 5704
rect 31300 5652 31352 5704
rect 31760 5652 31812 5704
rect 34612 5652 34664 5704
rect 35440 5652 35492 5704
rect 25872 5516 25924 5568
rect 27804 5516 27856 5568
rect 28540 5584 28592 5636
rect 29276 5584 29328 5636
rect 28724 5516 28776 5568
rect 29092 5559 29144 5568
rect 29092 5525 29101 5559
rect 29101 5525 29135 5559
rect 29135 5525 29144 5559
rect 29092 5516 29144 5525
rect 29184 5516 29236 5568
rect 30104 5559 30156 5568
rect 30104 5525 30113 5559
rect 30113 5525 30147 5559
rect 30147 5525 30156 5559
rect 30104 5516 30156 5525
rect 30380 5516 30432 5568
rect 30472 5516 30524 5568
rect 31208 5516 31260 5568
rect 32956 5584 33008 5636
rect 34244 5516 34296 5568
rect 35624 5516 35676 5568
rect 35900 5763 35952 5772
rect 35900 5729 35909 5763
rect 35909 5729 35943 5763
rect 35943 5729 35952 5763
rect 35900 5720 35952 5729
rect 36820 5720 36872 5772
rect 38016 5856 38068 5908
rect 37280 5652 37332 5704
rect 38384 5695 38436 5704
rect 38384 5661 38393 5695
rect 38393 5661 38427 5695
rect 38427 5661 38436 5695
rect 38384 5652 38436 5661
rect 36084 5584 36136 5636
rect 37188 5516 37240 5568
rect 10472 5414 10524 5466
rect 10536 5414 10588 5466
rect 10600 5414 10652 5466
rect 10664 5414 10716 5466
rect 10728 5414 10780 5466
rect 19994 5414 20046 5466
rect 20058 5414 20110 5466
rect 20122 5414 20174 5466
rect 20186 5414 20238 5466
rect 20250 5414 20302 5466
rect 29516 5414 29568 5466
rect 29580 5414 29632 5466
rect 29644 5414 29696 5466
rect 29708 5414 29760 5466
rect 29772 5414 29824 5466
rect 39038 5414 39090 5466
rect 39102 5414 39154 5466
rect 39166 5414 39218 5466
rect 39230 5414 39282 5466
rect 39294 5414 39346 5466
rect 1768 5355 1820 5364
rect 1768 5321 1777 5355
rect 1777 5321 1811 5355
rect 1811 5321 1820 5355
rect 1768 5312 1820 5321
rect 6092 5312 6144 5364
rect 2044 5244 2096 5296
rect 4344 5287 4396 5296
rect 4344 5253 4353 5287
rect 4353 5253 4387 5287
rect 4387 5253 4396 5287
rect 4344 5244 4396 5253
rect 6000 5287 6052 5296
rect 6000 5253 6009 5287
rect 6009 5253 6043 5287
rect 6043 5253 6052 5287
rect 6000 5244 6052 5253
rect 7288 5244 7340 5296
rect 9404 5312 9456 5364
rect 10968 5312 11020 5364
rect 15016 5312 15068 5364
rect 11060 5244 11112 5296
rect 11888 5244 11940 5296
rect 13268 5244 13320 5296
rect 13360 5244 13412 5296
rect 15476 5312 15528 5364
rect 15660 5312 15712 5364
rect 15292 5244 15344 5296
rect 940 5176 992 5228
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 8944 5176 8996 5228
rect 1584 5040 1636 5092
rect 2596 5151 2648 5160
rect 2596 5117 2605 5151
rect 2605 5117 2639 5151
rect 2639 5117 2648 5151
rect 2596 5108 2648 5117
rect 3884 5040 3936 5092
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 14096 5176 14148 5228
rect 17868 5312 17920 5364
rect 17960 5312 18012 5364
rect 17132 5287 17184 5296
rect 17132 5253 17141 5287
rect 17141 5253 17175 5287
rect 17175 5253 17184 5287
rect 17132 5244 17184 5253
rect 17592 5244 17644 5296
rect 18696 5244 18748 5296
rect 2412 4972 2464 5024
rect 10140 5108 10192 5160
rect 6920 4972 6972 5024
rect 7932 4972 7984 5024
rect 8208 4972 8260 5024
rect 9036 4972 9088 5024
rect 9496 4972 9548 5024
rect 11336 5108 11388 5160
rect 11980 5151 12032 5160
rect 11980 5117 11989 5151
rect 11989 5117 12023 5151
rect 12023 5117 12032 5151
rect 11980 5108 12032 5117
rect 13912 4972 13964 5024
rect 14832 5151 14884 5160
rect 14832 5117 14841 5151
rect 14841 5117 14875 5151
rect 14875 5117 14884 5151
rect 14832 5108 14884 5117
rect 15384 5108 15436 5160
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 16120 5040 16172 5092
rect 20812 5312 20864 5364
rect 21364 5287 21416 5296
rect 21364 5253 21373 5287
rect 21373 5253 21407 5287
rect 21407 5253 21416 5287
rect 21364 5244 21416 5253
rect 21640 5244 21692 5296
rect 22376 5244 22428 5296
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 22468 5176 22520 5228
rect 22284 5108 22336 5160
rect 23020 5244 23072 5296
rect 22928 5176 22980 5228
rect 14924 4972 14976 5024
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16304 4972 16356 4981
rect 20352 5040 20404 5092
rect 23848 5151 23900 5160
rect 23848 5117 23857 5151
rect 23857 5117 23891 5151
rect 23891 5117 23900 5151
rect 23848 5108 23900 5117
rect 24676 5176 24728 5228
rect 25136 5244 25188 5296
rect 26884 5244 26936 5296
rect 27344 5287 27396 5296
rect 27344 5253 27353 5287
rect 27353 5253 27387 5287
rect 27387 5253 27396 5287
rect 27344 5244 27396 5253
rect 28172 5312 28224 5364
rect 29368 5312 29420 5364
rect 30288 5312 30340 5364
rect 32128 5312 32180 5364
rect 34704 5312 34756 5364
rect 34796 5312 34848 5364
rect 35716 5312 35768 5364
rect 28540 5244 28592 5296
rect 29920 5244 29972 5296
rect 24032 5108 24084 5160
rect 19064 4972 19116 5024
rect 19432 4972 19484 5024
rect 24032 4972 24084 5024
rect 26976 5108 27028 5160
rect 27528 5219 27580 5228
rect 27528 5185 27537 5219
rect 27537 5185 27571 5219
rect 27571 5185 27580 5219
rect 27528 5176 27580 5185
rect 28172 5219 28224 5228
rect 28172 5185 28181 5219
rect 28181 5185 28215 5219
rect 28215 5185 28224 5219
rect 28172 5176 28224 5185
rect 28080 5040 28132 5092
rect 27344 4972 27396 5024
rect 29184 5108 29236 5160
rect 30564 5176 30616 5228
rect 30840 5219 30892 5228
rect 30840 5185 30849 5219
rect 30849 5185 30883 5219
rect 30883 5185 30892 5219
rect 30840 5176 30892 5185
rect 31300 5176 31352 5228
rect 32128 5176 32180 5228
rect 32404 5219 32456 5228
rect 32404 5185 32413 5219
rect 32413 5185 32447 5219
rect 32447 5185 32456 5219
rect 32404 5176 32456 5185
rect 33508 5244 33560 5296
rect 36636 5312 36688 5364
rect 36912 5312 36964 5364
rect 37464 5312 37516 5364
rect 37832 5244 37884 5296
rect 35256 5176 35308 5228
rect 35716 5219 35768 5228
rect 35716 5185 35725 5219
rect 35725 5185 35759 5219
rect 35759 5185 35768 5219
rect 35716 5176 35768 5185
rect 30932 5151 30984 5160
rect 30932 5117 30941 5151
rect 30941 5117 30975 5151
rect 30975 5117 30984 5151
rect 30932 5108 30984 5117
rect 33416 5151 33468 5160
rect 33416 5117 33425 5151
rect 33425 5117 33459 5151
rect 33459 5117 33468 5151
rect 33416 5108 33468 5117
rect 33876 5108 33928 5160
rect 35992 5176 36044 5228
rect 37464 5219 37516 5228
rect 37464 5185 37473 5219
rect 37473 5185 37507 5219
rect 37507 5185 37516 5219
rect 37464 5176 37516 5185
rect 38108 5219 38160 5228
rect 38108 5185 38117 5219
rect 38117 5185 38151 5219
rect 38151 5185 38160 5219
rect 38108 5176 38160 5185
rect 33048 5040 33100 5092
rect 30104 4972 30156 5024
rect 30380 5015 30432 5024
rect 30380 4981 30389 5015
rect 30389 4981 30423 5015
rect 30423 4981 30432 5015
rect 30380 4972 30432 4981
rect 31944 4972 31996 5024
rect 36912 5083 36964 5092
rect 36912 5049 36921 5083
rect 36921 5049 36955 5083
rect 36955 5049 36964 5083
rect 36912 5040 36964 5049
rect 34704 4972 34756 5024
rect 35992 4972 36044 5024
rect 36728 5015 36780 5024
rect 36728 4981 36737 5015
rect 36737 4981 36771 5015
rect 36771 4981 36780 5015
rect 36728 4972 36780 4981
rect 5711 4870 5763 4922
rect 5775 4870 5827 4922
rect 5839 4870 5891 4922
rect 5903 4870 5955 4922
rect 5967 4870 6019 4922
rect 15233 4870 15285 4922
rect 15297 4870 15349 4922
rect 15361 4870 15413 4922
rect 15425 4870 15477 4922
rect 15489 4870 15541 4922
rect 24755 4870 24807 4922
rect 24819 4870 24871 4922
rect 24883 4870 24935 4922
rect 24947 4870 24999 4922
rect 25011 4870 25063 4922
rect 34277 4870 34329 4922
rect 34341 4870 34393 4922
rect 34405 4870 34457 4922
rect 34469 4870 34521 4922
rect 34533 4870 34585 4922
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 4896 4768 4948 4820
rect 5080 4768 5132 4820
rect 8576 4768 8628 4820
rect 9220 4768 9272 4820
rect 11060 4768 11112 4820
rect 11980 4768 12032 4820
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 3332 4675 3384 4684
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 6092 4700 6144 4752
rect 8208 4700 8260 4752
rect 3332 4632 3384 4641
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 3700 4564 3752 4616
rect 2504 4496 2556 4548
rect 5172 4632 5224 4684
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 6552 4632 6604 4684
rect 6828 4632 6880 4684
rect 9772 4632 9824 4684
rect 17132 4768 17184 4820
rect 17592 4768 17644 4820
rect 21272 4768 21324 4820
rect 22008 4768 22060 4820
rect 14188 4700 14240 4752
rect 10876 4675 10928 4684
rect 10876 4641 10885 4675
rect 10885 4641 10919 4675
rect 10919 4641 10928 4675
rect 10876 4632 10928 4641
rect 10968 4632 11020 4684
rect 12256 4632 12308 4684
rect 12440 4632 12492 4684
rect 13360 4632 13412 4684
rect 13452 4675 13504 4684
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 14740 4700 14792 4752
rect 16580 4700 16632 4752
rect 13452 4632 13504 4641
rect 14556 4632 14608 4684
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 5908 4564 5960 4616
rect 8300 4564 8352 4616
rect 8576 4564 8628 4616
rect 4620 4428 4672 4480
rect 5080 4428 5132 4480
rect 5172 4428 5224 4480
rect 5724 4496 5776 4548
rect 7748 4496 7800 4548
rect 7932 4428 7984 4480
rect 9680 4564 9732 4616
rect 9220 4539 9272 4548
rect 9220 4505 9229 4539
rect 9229 4505 9263 4539
rect 9263 4505 9272 4539
rect 9220 4496 9272 4505
rect 11152 4564 11204 4616
rect 11244 4564 11296 4616
rect 12992 4564 13044 4616
rect 13912 4564 13964 4616
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14924 4632 14976 4684
rect 15660 4632 15712 4684
rect 17684 4632 17736 4684
rect 18328 4632 18380 4684
rect 20536 4700 20588 4752
rect 22192 4700 22244 4752
rect 22928 4700 22980 4752
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 19984 4675 20036 4684
rect 19984 4641 19993 4675
rect 19993 4641 20027 4675
rect 20027 4641 20036 4675
rect 19984 4632 20036 4641
rect 22652 4632 22704 4684
rect 14556 4539 14608 4548
rect 14556 4505 14565 4539
rect 14565 4505 14599 4539
rect 14599 4505 14608 4539
rect 14556 4496 14608 4505
rect 16672 4564 16724 4616
rect 16948 4564 17000 4616
rect 15476 4496 15528 4548
rect 15568 4539 15620 4548
rect 15568 4505 15577 4539
rect 15577 4505 15611 4539
rect 15611 4505 15620 4539
rect 15568 4496 15620 4505
rect 9680 4428 9732 4480
rect 12164 4428 12216 4480
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 14280 4428 14332 4480
rect 19248 4496 19300 4548
rect 19432 4564 19484 4616
rect 20628 4607 20680 4616
rect 20628 4573 20637 4607
rect 20637 4573 20671 4607
rect 20671 4573 20680 4607
rect 20628 4564 20680 4573
rect 22836 4564 22888 4616
rect 23204 4607 23256 4616
rect 23204 4573 23213 4607
rect 23213 4573 23247 4607
rect 23247 4573 23256 4607
rect 23204 4564 23256 4573
rect 23940 4700 23992 4752
rect 25780 4811 25832 4820
rect 25780 4777 25789 4811
rect 25789 4777 25823 4811
rect 25823 4777 25832 4811
rect 25780 4768 25832 4777
rect 26056 4811 26108 4820
rect 26056 4777 26065 4811
rect 26065 4777 26099 4811
rect 26099 4777 26108 4811
rect 26056 4768 26108 4777
rect 23388 4632 23440 4684
rect 23572 4607 23624 4616
rect 23572 4573 23581 4607
rect 23581 4573 23615 4607
rect 23615 4573 23624 4607
rect 23572 4564 23624 4573
rect 24400 4564 24452 4616
rect 26332 4607 26384 4616
rect 26332 4573 26341 4607
rect 26341 4573 26375 4607
rect 26375 4573 26384 4607
rect 26332 4564 26384 4573
rect 27436 4768 27488 4820
rect 29000 4768 29052 4820
rect 30104 4768 30156 4820
rect 34428 4768 34480 4820
rect 36176 4768 36228 4820
rect 36544 4768 36596 4820
rect 37188 4768 37240 4820
rect 27252 4632 27304 4684
rect 29000 4632 29052 4684
rect 28172 4607 28224 4616
rect 28172 4573 28181 4607
rect 28181 4573 28215 4607
rect 28215 4573 28224 4607
rect 28172 4564 28224 4573
rect 28356 4607 28408 4616
rect 28356 4573 28365 4607
rect 28365 4573 28399 4607
rect 28399 4573 28408 4607
rect 28356 4564 28408 4573
rect 28540 4607 28592 4616
rect 28540 4573 28549 4607
rect 28549 4573 28583 4607
rect 28583 4573 28592 4607
rect 28540 4564 28592 4573
rect 23480 4496 23532 4548
rect 23848 4496 23900 4548
rect 24768 4496 24820 4548
rect 18512 4471 18564 4480
rect 18512 4437 18521 4471
rect 18521 4437 18555 4471
rect 18555 4437 18564 4471
rect 18512 4428 18564 4437
rect 19616 4428 19668 4480
rect 20260 4428 20312 4480
rect 21272 4428 21324 4480
rect 25780 4496 25832 4548
rect 26240 4496 26292 4548
rect 28264 4496 28316 4548
rect 28448 4539 28500 4548
rect 28448 4505 28457 4539
rect 28457 4505 28491 4539
rect 28491 4505 28500 4539
rect 28448 4496 28500 4505
rect 27528 4428 27580 4480
rect 31024 4700 31076 4752
rect 30012 4675 30064 4684
rect 30012 4641 30021 4675
rect 30021 4641 30055 4675
rect 30055 4641 30064 4675
rect 30012 4632 30064 4641
rect 32036 4675 32088 4684
rect 32036 4641 32045 4675
rect 32045 4641 32079 4675
rect 32079 4641 32088 4675
rect 32036 4632 32088 4641
rect 33048 4632 33100 4684
rect 29368 4564 29420 4616
rect 31944 4564 31996 4616
rect 35072 4564 35124 4616
rect 36176 4564 36228 4616
rect 30012 4496 30064 4548
rect 30288 4496 30340 4548
rect 33784 4496 33836 4548
rect 37188 4607 37240 4616
rect 37188 4573 37197 4607
rect 37197 4573 37231 4607
rect 37231 4573 37240 4607
rect 37188 4564 37240 4573
rect 37096 4496 37148 4548
rect 37556 4564 37608 4616
rect 37464 4496 37516 4548
rect 38384 4496 38436 4548
rect 32128 4428 32180 4480
rect 34428 4428 34480 4480
rect 34796 4428 34848 4480
rect 38292 4428 38344 4480
rect 10472 4326 10524 4378
rect 10536 4326 10588 4378
rect 10600 4326 10652 4378
rect 10664 4326 10716 4378
rect 10728 4326 10780 4378
rect 19994 4326 20046 4378
rect 20058 4326 20110 4378
rect 20122 4326 20174 4378
rect 20186 4326 20238 4378
rect 20250 4326 20302 4378
rect 29516 4326 29568 4378
rect 29580 4326 29632 4378
rect 29644 4326 29696 4378
rect 29708 4326 29760 4378
rect 29772 4326 29824 4378
rect 39038 4326 39090 4378
rect 39102 4326 39154 4378
rect 39166 4326 39218 4378
rect 39230 4326 39282 4378
rect 39294 4326 39346 4378
rect 5448 4224 5500 4276
rect 2964 4156 3016 4208
rect 5172 4156 5224 4208
rect 8484 4224 8536 4276
rect 13360 4224 13412 4276
rect 13912 4224 13964 4276
rect 14004 4224 14056 4276
rect 5908 4156 5960 4208
rect 1584 4020 1636 4072
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 3424 4020 3476 4072
rect 5632 4088 5684 4140
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 7288 4156 7340 4208
rect 8208 4156 8260 4208
rect 10324 4156 10376 4208
rect 10692 4199 10744 4208
rect 10692 4165 10701 4199
rect 10701 4165 10735 4199
rect 10735 4165 10744 4199
rect 10692 4156 10744 4165
rect 13452 4156 13504 4208
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 5816 4020 5868 4072
rect 5908 4063 5960 4072
rect 5908 4029 5917 4063
rect 5917 4029 5951 4063
rect 5951 4029 5960 4063
rect 5908 4020 5960 4029
rect 6552 4020 6604 4072
rect 7104 4088 7156 4140
rect 7932 4088 7984 4140
rect 8116 4063 8168 4072
rect 4344 3952 4396 4004
rect 1768 3927 1820 3936
rect 1768 3893 1777 3927
rect 1777 3893 1811 3927
rect 1811 3893 1820 3927
rect 1768 3884 1820 3893
rect 5356 3884 5408 3936
rect 5632 3884 5684 3936
rect 6736 3884 6788 3936
rect 7012 3952 7064 4004
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 14832 4156 14884 4208
rect 15200 4156 15252 4208
rect 10232 4088 10284 4140
rect 9680 4020 9732 4072
rect 10140 4020 10192 4072
rect 12072 4088 12124 4140
rect 12348 4131 12400 4140
rect 12348 4097 12357 4131
rect 12357 4097 12391 4131
rect 12391 4097 12400 4131
rect 12348 4088 12400 4097
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 12992 4020 13044 4072
rect 14280 4131 14332 4140
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 14188 4020 14240 4072
rect 14648 4020 14700 4072
rect 15568 4020 15620 4072
rect 17592 4156 17644 4208
rect 20444 4224 20496 4276
rect 19524 4156 19576 4208
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 17040 4088 17092 4140
rect 17224 4131 17276 4140
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 17316 4131 17368 4140
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 17868 4088 17920 4140
rect 20996 4156 21048 4208
rect 22284 4224 22336 4276
rect 22928 4224 22980 4276
rect 24492 4224 24544 4276
rect 26240 4224 26292 4276
rect 28172 4224 28224 4276
rect 31944 4224 31996 4276
rect 21640 4088 21692 4140
rect 24032 4088 24084 4140
rect 24860 4131 24912 4140
rect 24860 4097 24869 4131
rect 24869 4097 24903 4131
rect 24903 4097 24912 4131
rect 24860 4088 24912 4097
rect 26608 4156 26660 4208
rect 28080 4156 28132 4208
rect 7656 3927 7708 3936
rect 7656 3893 7665 3927
rect 7665 3893 7699 3927
rect 7699 3893 7708 3927
rect 7656 3884 7708 3893
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10140 3884 10192 3893
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 12808 3952 12860 4004
rect 13912 3952 13964 4004
rect 13636 3884 13688 3936
rect 14096 3884 14148 3936
rect 17776 4020 17828 4072
rect 17132 3952 17184 4004
rect 20352 4020 20404 4072
rect 21364 4063 21416 4072
rect 21364 4029 21373 4063
rect 21373 4029 21407 4063
rect 21407 4029 21416 4063
rect 21364 4020 21416 4029
rect 19340 3952 19392 4004
rect 20628 3952 20680 4004
rect 22560 4063 22612 4072
rect 22560 4029 22569 4063
rect 22569 4029 22603 4063
rect 22603 4029 22612 4063
rect 22560 4020 22612 4029
rect 22652 4020 22704 4072
rect 15752 3884 15804 3936
rect 17316 3884 17368 3936
rect 19524 3884 19576 3936
rect 22192 3884 22244 3936
rect 24676 3952 24728 4004
rect 25136 4063 25188 4072
rect 25136 4029 25145 4063
rect 25145 4029 25179 4063
rect 25179 4029 25188 4063
rect 25136 4020 25188 4029
rect 26240 4063 26292 4072
rect 26240 4029 26249 4063
rect 26249 4029 26283 4063
rect 26283 4029 26292 4063
rect 26240 4020 26292 4029
rect 24492 3927 24544 3936
rect 24492 3893 24501 3927
rect 24501 3893 24535 3927
rect 24535 3893 24544 3927
rect 24492 3884 24544 3893
rect 25688 3927 25740 3936
rect 25688 3893 25697 3927
rect 25697 3893 25731 3927
rect 25731 3893 25740 3927
rect 25688 3884 25740 3893
rect 27252 3884 27304 3936
rect 27712 3884 27764 3936
rect 28264 3952 28316 4004
rect 28724 4088 28776 4140
rect 28632 4063 28684 4072
rect 28632 4029 28641 4063
rect 28641 4029 28675 4063
rect 28675 4029 28684 4063
rect 28632 4020 28684 4029
rect 30012 4156 30064 4208
rect 35164 4224 35216 4276
rect 35808 4224 35860 4276
rect 35992 4224 36044 4276
rect 33600 4156 33652 4208
rect 35440 4199 35492 4208
rect 35440 4165 35449 4199
rect 35449 4165 35483 4199
rect 35483 4165 35492 4199
rect 35440 4156 35492 4165
rect 35624 4156 35676 4208
rect 32036 4088 32088 4140
rect 37280 4088 37332 4140
rect 38108 4131 38160 4140
rect 38108 4097 38117 4131
rect 38117 4097 38151 4131
rect 38151 4097 38160 4131
rect 38108 4088 38160 4097
rect 29460 4063 29512 4072
rect 29460 4029 29469 4063
rect 29469 4029 29503 4063
rect 29503 4029 29512 4063
rect 29460 4020 29512 4029
rect 30380 4020 30432 4072
rect 32680 4020 32732 4072
rect 32956 4020 33008 4072
rect 32128 3952 32180 4004
rect 34980 4020 35032 4072
rect 30840 3884 30892 3936
rect 33140 3884 33192 3936
rect 36084 3884 36136 3936
rect 36268 3952 36320 4004
rect 38200 3927 38252 3936
rect 38200 3893 38209 3927
rect 38209 3893 38243 3927
rect 38243 3893 38252 3927
rect 38200 3884 38252 3893
rect 5711 3782 5763 3834
rect 5775 3782 5827 3834
rect 5839 3782 5891 3834
rect 5903 3782 5955 3834
rect 5967 3782 6019 3834
rect 15233 3782 15285 3834
rect 15297 3782 15349 3834
rect 15361 3782 15413 3834
rect 15425 3782 15477 3834
rect 15489 3782 15541 3834
rect 24755 3782 24807 3834
rect 24819 3782 24871 3834
rect 24883 3782 24935 3834
rect 24947 3782 24999 3834
rect 25011 3782 25063 3834
rect 34277 3782 34329 3834
rect 34341 3782 34393 3834
rect 34405 3782 34457 3834
rect 34469 3782 34521 3834
rect 34533 3782 34585 3834
rect 2596 3680 2648 3732
rect 3976 3723 4028 3732
rect 3976 3689 3985 3723
rect 3985 3689 4019 3723
rect 4019 3689 4028 3723
rect 3976 3680 4028 3689
rect 8208 3680 8260 3732
rect 12164 3680 12216 3732
rect 1676 3612 1728 3664
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 3516 3544 3568 3596
rect 4436 3544 4488 3596
rect 1308 3476 1360 3528
rect 2780 3476 2832 3528
rect 4252 3476 4304 3528
rect 4620 3476 4672 3528
rect 6276 3612 6328 3664
rect 6552 3612 6604 3664
rect 14648 3612 14700 3664
rect 16304 3680 16356 3732
rect 18512 3680 18564 3732
rect 18604 3680 18656 3732
rect 5632 3544 5684 3596
rect 6000 3587 6052 3596
rect 6000 3553 6009 3587
rect 6009 3553 6043 3587
rect 6043 3553 6052 3587
rect 6000 3544 6052 3553
rect 6736 3544 6788 3596
rect 7104 3544 7156 3596
rect 7288 3587 7340 3596
rect 7288 3553 7297 3587
rect 7297 3553 7331 3587
rect 7331 3553 7340 3587
rect 7288 3544 7340 3553
rect 8760 3544 8812 3596
rect 10048 3587 10100 3596
rect 10048 3553 10057 3587
rect 10057 3553 10091 3587
rect 10091 3553 10100 3587
rect 10048 3544 10100 3553
rect 10140 3544 10192 3596
rect 12348 3544 12400 3596
rect 14924 3587 14976 3596
rect 14924 3553 14933 3587
rect 14933 3553 14967 3587
rect 14967 3553 14976 3587
rect 14924 3544 14976 3553
rect 16580 3544 16632 3596
rect 8392 3476 8444 3528
rect 11060 3476 11112 3528
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 12992 3476 13044 3528
rect 13820 3476 13872 3528
rect 14096 3476 14148 3528
rect 16856 3544 16908 3596
rect 17132 3587 17184 3596
rect 17132 3553 17141 3587
rect 17141 3553 17175 3587
rect 17175 3553 17184 3587
rect 17132 3544 17184 3553
rect 17776 3544 17828 3596
rect 19892 3680 19944 3732
rect 19432 3587 19484 3596
rect 19432 3553 19441 3587
rect 19441 3553 19475 3587
rect 19475 3553 19484 3587
rect 19432 3544 19484 3553
rect 22560 3680 22612 3732
rect 25688 3680 25740 3732
rect 27344 3680 27396 3732
rect 27436 3723 27488 3732
rect 27436 3689 27445 3723
rect 27445 3689 27479 3723
rect 27479 3689 27488 3723
rect 27436 3680 27488 3689
rect 28356 3680 28408 3732
rect 28908 3680 28960 3732
rect 29000 3680 29052 3732
rect 33048 3680 33100 3732
rect 37280 3680 37332 3732
rect 22652 3544 22704 3596
rect 22928 3587 22980 3596
rect 22928 3553 22937 3587
rect 22937 3553 22971 3587
rect 22971 3553 22980 3587
rect 22928 3544 22980 3553
rect 23204 3544 23256 3596
rect 2872 3408 2924 3460
rect 9680 3408 9732 3460
rect 11612 3451 11664 3460
rect 11612 3417 11621 3451
rect 11621 3417 11655 3451
rect 11655 3417 11664 3451
rect 11612 3408 11664 3417
rect 12624 3408 12676 3460
rect 5172 3340 5224 3392
rect 6368 3340 6420 3392
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 15476 3408 15528 3460
rect 16488 3408 16540 3460
rect 7104 3340 7156 3349
rect 13084 3383 13136 3392
rect 13084 3349 13093 3383
rect 13093 3349 13127 3383
rect 13127 3349 13136 3383
rect 13084 3340 13136 3349
rect 16948 3340 17000 3392
rect 20812 3476 20864 3528
rect 17408 3451 17460 3460
rect 17408 3417 17417 3451
rect 17417 3417 17451 3451
rect 17451 3417 17460 3451
rect 17408 3408 17460 3417
rect 17960 3408 18012 3460
rect 19800 3408 19852 3460
rect 19524 3340 19576 3392
rect 23388 3476 23440 3528
rect 24400 3544 24452 3596
rect 24676 3544 24728 3596
rect 31944 3612 31996 3664
rect 21088 3408 21140 3460
rect 24032 3476 24084 3528
rect 26148 3476 26200 3528
rect 27252 3519 27304 3528
rect 27252 3485 27261 3519
rect 27261 3485 27295 3519
rect 27295 3485 27304 3519
rect 27252 3476 27304 3485
rect 21272 3340 21324 3392
rect 26608 3408 26660 3460
rect 27528 3408 27580 3460
rect 28448 3451 28500 3460
rect 28448 3417 28457 3451
rect 28457 3417 28491 3451
rect 28491 3417 28500 3451
rect 28448 3408 28500 3417
rect 29460 3544 29512 3596
rect 32036 3544 32088 3596
rect 28908 3476 28960 3528
rect 29644 3476 29696 3528
rect 30104 3476 30156 3528
rect 36636 3655 36688 3664
rect 36636 3621 36645 3655
rect 36645 3621 36679 3655
rect 36679 3621 36688 3655
rect 36636 3612 36688 3621
rect 32404 3544 32456 3596
rect 34888 3587 34940 3596
rect 34888 3553 34897 3587
rect 34897 3553 34931 3587
rect 34931 3553 34940 3587
rect 34888 3544 34940 3553
rect 35808 3544 35860 3596
rect 37004 3544 37056 3596
rect 34060 3476 34112 3528
rect 37096 3476 37148 3528
rect 28264 3340 28316 3392
rect 30472 3408 30524 3460
rect 34796 3408 34848 3460
rect 35164 3451 35216 3460
rect 35164 3417 35173 3451
rect 35173 3417 35207 3451
rect 35207 3417 35216 3451
rect 35164 3408 35216 3417
rect 31484 3340 31536 3392
rect 33324 3340 33376 3392
rect 33600 3340 33652 3392
rect 35900 3340 35952 3392
rect 38660 3451 38712 3460
rect 38660 3417 38669 3451
rect 38669 3417 38703 3451
rect 38703 3417 38712 3451
rect 38660 3408 38712 3417
rect 37280 3383 37332 3392
rect 37280 3349 37289 3383
rect 37289 3349 37323 3383
rect 37323 3349 37332 3383
rect 37280 3340 37332 3349
rect 10472 3238 10524 3290
rect 10536 3238 10588 3290
rect 10600 3238 10652 3290
rect 10664 3238 10716 3290
rect 10728 3238 10780 3290
rect 19994 3238 20046 3290
rect 20058 3238 20110 3290
rect 20122 3238 20174 3290
rect 20186 3238 20238 3290
rect 20250 3238 20302 3290
rect 29516 3238 29568 3290
rect 29580 3238 29632 3290
rect 29644 3238 29696 3290
rect 29708 3238 29760 3290
rect 29772 3238 29824 3290
rect 39038 3238 39090 3290
rect 39102 3238 39154 3290
rect 39166 3238 39218 3290
rect 39230 3238 39282 3290
rect 39294 3238 39346 3290
rect 5264 3136 5316 3188
rect 5724 3179 5776 3188
rect 5724 3145 5733 3179
rect 5733 3145 5767 3179
rect 5767 3145 5776 3179
rect 5724 3136 5776 3145
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 7288 3136 7340 3188
rect 8116 3136 8168 3188
rect 11612 3136 11664 3188
rect 12164 3179 12216 3188
rect 12164 3145 12173 3179
rect 12173 3145 12207 3179
rect 12207 3145 12216 3179
rect 12164 3136 12216 3145
rect 13084 3136 13136 3188
rect 13360 3136 13412 3188
rect 15476 3136 15528 3188
rect 1860 3111 1912 3120
rect 1860 3077 1869 3111
rect 1869 3077 1903 3111
rect 1903 3077 1912 3111
rect 1860 3068 1912 3077
rect 3424 3068 3476 3120
rect 4160 3068 4212 3120
rect 6092 3068 6144 3120
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 3792 3000 3844 3052
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 4804 3000 4856 3052
rect 3700 2932 3752 2984
rect 5724 3000 5776 3052
rect 7656 3068 7708 3120
rect 9864 3068 9916 3120
rect 11244 3068 11296 3120
rect 11336 3068 11388 3120
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 7564 3000 7616 3052
rect 8208 3000 8260 3052
rect 6092 2932 6144 2984
rect 7012 2932 7064 2984
rect 7932 2975 7984 2984
rect 7932 2941 7941 2975
rect 7941 2941 7975 2975
rect 7975 2941 7984 2975
rect 7932 2932 7984 2941
rect 6828 2864 6880 2916
rect 8852 2932 8904 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 14188 3068 14240 3120
rect 14372 3068 14424 3120
rect 19892 3136 19944 3188
rect 27068 3136 27120 3188
rect 27252 3136 27304 3188
rect 19616 3111 19668 3120
rect 19616 3077 19625 3111
rect 19625 3077 19659 3111
rect 19659 3077 19668 3111
rect 19616 3068 19668 3077
rect 20904 3068 20956 3120
rect 22192 3068 22244 3120
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 18236 3000 18288 3052
rect 19340 3043 19392 3052
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 23388 3000 23440 3052
rect 24584 3068 24636 3120
rect 26056 3068 26108 3120
rect 27896 3068 27948 3120
rect 25780 3000 25832 3052
rect 27344 3000 27396 3052
rect 27528 3043 27580 3052
rect 27528 3009 27537 3043
rect 27537 3009 27571 3043
rect 27571 3009 27580 3043
rect 27528 3000 27580 3009
rect 29000 3068 29052 3120
rect 32128 3136 32180 3188
rect 16764 2932 16816 2984
rect 22008 2975 22060 2984
rect 22008 2941 22017 2975
rect 22017 2941 22051 2975
rect 22051 2941 22060 2975
rect 22008 2932 22060 2941
rect 11152 2907 11204 2916
rect 11152 2873 11161 2907
rect 11161 2873 11195 2907
rect 11195 2873 11204 2907
rect 11152 2864 11204 2873
rect 22744 2932 22796 2984
rect 24124 2932 24176 2984
rect 24860 2932 24912 2984
rect 28080 3000 28132 3052
rect 28540 2932 28592 2984
rect 30012 3000 30064 3052
rect 28908 2975 28960 2984
rect 28908 2941 28917 2975
rect 28917 2941 28951 2975
rect 28951 2941 28960 2975
rect 28908 2932 28960 2941
rect 6736 2796 6788 2848
rect 6920 2796 6972 2848
rect 11060 2796 11112 2848
rect 14004 2796 14056 2848
rect 14096 2796 14148 2848
rect 19340 2796 19392 2848
rect 25504 2864 25556 2916
rect 20904 2796 20956 2848
rect 24308 2796 24360 2848
rect 27620 2796 27672 2848
rect 28080 2796 28132 2848
rect 31852 3000 31904 3052
rect 32496 3111 32548 3120
rect 32496 3077 32505 3111
rect 32505 3077 32539 3111
rect 32539 3077 32548 3111
rect 32496 3068 32548 3077
rect 33968 3136 34020 3188
rect 33416 3111 33468 3120
rect 33416 3077 33425 3111
rect 33425 3077 33459 3111
rect 33459 3077 33468 3111
rect 33416 3068 33468 3077
rect 37464 3136 37516 3188
rect 34704 3068 34756 3120
rect 36820 3068 36872 3120
rect 34888 3000 34940 3052
rect 37096 3000 37148 3052
rect 30104 2796 30156 2848
rect 30380 2839 30432 2848
rect 30380 2805 30389 2839
rect 30389 2805 30423 2839
rect 30423 2805 30432 2839
rect 30380 2796 30432 2805
rect 33508 2932 33560 2984
rect 32312 2864 32364 2916
rect 36820 2975 36872 2984
rect 36820 2941 36829 2975
rect 36829 2941 36863 2975
rect 36863 2941 36872 2975
rect 36820 2932 36872 2941
rect 39396 2864 39448 2916
rect 33048 2796 33100 2848
rect 33140 2796 33192 2848
rect 37556 2839 37608 2848
rect 37556 2805 37565 2839
rect 37565 2805 37599 2839
rect 37599 2805 37608 2839
rect 37556 2796 37608 2805
rect 5711 2694 5763 2746
rect 5775 2694 5827 2746
rect 5839 2694 5891 2746
rect 5903 2694 5955 2746
rect 5967 2694 6019 2746
rect 15233 2694 15285 2746
rect 15297 2694 15349 2746
rect 15361 2694 15413 2746
rect 15425 2694 15477 2746
rect 15489 2694 15541 2746
rect 24755 2694 24807 2746
rect 24819 2694 24871 2746
rect 24883 2694 24935 2746
rect 24947 2694 24999 2746
rect 25011 2694 25063 2746
rect 34277 2694 34329 2746
rect 34341 2694 34393 2746
rect 34405 2694 34457 2746
rect 34469 2694 34521 2746
rect 34533 2694 34585 2746
rect 4712 2592 4764 2644
rect 12900 2592 12952 2644
rect 7840 2524 7892 2576
rect 9496 2524 9548 2576
rect 3608 2456 3660 2508
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 5632 2456 5684 2508
rect 4804 2431 4856 2440
rect 4804 2397 4813 2431
rect 4813 2397 4847 2431
rect 4847 2397 4856 2431
rect 4804 2388 4856 2397
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6460 2456 6512 2508
rect 6828 2456 6880 2508
rect 8392 2456 8444 2508
rect 11796 2567 11848 2576
rect 11796 2533 11805 2567
rect 11805 2533 11839 2567
rect 11839 2533 11848 2567
rect 11796 2524 11848 2533
rect 11888 2524 11940 2576
rect 12992 2524 13044 2576
rect 15844 2592 15896 2644
rect 17868 2592 17920 2644
rect 18144 2592 18196 2644
rect 21180 2635 21232 2644
rect 21180 2601 21189 2635
rect 21189 2601 21223 2635
rect 21223 2601 21232 2635
rect 21180 2592 21232 2601
rect 24492 2592 24544 2644
rect 26332 2635 26384 2644
rect 26332 2601 26341 2635
rect 26341 2601 26375 2635
rect 26375 2601 26384 2635
rect 26332 2592 26384 2601
rect 26884 2592 26936 2644
rect 23848 2524 23900 2576
rect 28724 2592 28776 2644
rect 30656 2592 30708 2644
rect 33692 2592 33744 2644
rect 35532 2524 35584 2576
rect 3240 2363 3292 2372
rect 3240 2329 3249 2363
rect 3249 2329 3283 2363
rect 3283 2329 3292 2363
rect 3240 2320 3292 2329
rect 4160 2320 4212 2372
rect 4712 2363 4764 2372
rect 4712 2329 4721 2363
rect 4721 2329 4755 2363
rect 4755 2329 4764 2363
rect 4712 2320 4764 2329
rect 6184 2388 6236 2440
rect 8576 2388 8628 2440
rect 5540 2252 5592 2304
rect 6736 2320 6788 2372
rect 8944 2320 8996 2372
rect 10048 2388 10100 2440
rect 11888 2388 11940 2440
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 16856 2499 16908 2508
rect 16856 2465 16865 2499
rect 16865 2465 16899 2499
rect 16899 2465 16908 2499
rect 16856 2456 16908 2465
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 17224 2456 17276 2508
rect 17500 2456 17552 2508
rect 22008 2456 22060 2508
rect 24584 2499 24636 2508
rect 24584 2465 24593 2499
rect 24593 2465 24627 2499
rect 24627 2465 24636 2499
rect 24584 2456 24636 2465
rect 27528 2456 27580 2508
rect 31300 2456 31352 2508
rect 8484 2252 8536 2304
rect 12072 2363 12124 2372
rect 12072 2329 12081 2363
rect 12081 2329 12115 2363
rect 12115 2329 12124 2363
rect 12072 2320 12124 2329
rect 12164 2252 12216 2304
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 30104 2388 30156 2440
rect 30196 2388 30248 2440
rect 13176 2320 13228 2372
rect 14556 2363 14608 2372
rect 14556 2329 14565 2363
rect 14565 2329 14599 2363
rect 14599 2329 14608 2363
rect 14556 2320 14608 2329
rect 15200 2320 15252 2372
rect 18420 2320 18472 2372
rect 21088 2363 21140 2372
rect 21088 2329 21097 2363
rect 21097 2329 21131 2363
rect 21131 2329 21140 2363
rect 21088 2320 21140 2329
rect 24584 2320 24636 2372
rect 25136 2320 25188 2372
rect 25320 2320 25372 2372
rect 27712 2320 27764 2372
rect 29920 2320 29972 2372
rect 30748 2363 30800 2372
rect 30748 2329 30757 2363
rect 30757 2329 30791 2363
rect 30791 2329 30800 2363
rect 30748 2320 30800 2329
rect 32036 2456 32088 2508
rect 32588 2456 32640 2508
rect 34060 2388 34112 2440
rect 35440 2388 35492 2440
rect 17224 2252 17276 2304
rect 17868 2252 17920 2304
rect 27252 2252 27304 2304
rect 27344 2252 27396 2304
rect 29276 2252 29328 2304
rect 31668 2295 31720 2304
rect 31668 2261 31677 2295
rect 31677 2261 31711 2295
rect 31711 2261 31720 2295
rect 31668 2252 31720 2261
rect 33232 2320 33284 2372
rect 34152 2320 34204 2372
rect 35716 2320 35768 2372
rect 38476 2363 38528 2372
rect 38476 2329 38485 2363
rect 38485 2329 38519 2363
rect 38519 2329 38528 2363
rect 38476 2320 38528 2329
rect 38660 2363 38712 2372
rect 38660 2329 38669 2363
rect 38669 2329 38703 2363
rect 38703 2329 38712 2363
rect 38660 2320 38712 2329
rect 34060 2252 34112 2304
rect 36636 2295 36688 2304
rect 36636 2261 36645 2295
rect 36645 2261 36679 2295
rect 36679 2261 36688 2295
rect 36636 2252 36688 2261
rect 37648 2295 37700 2304
rect 37648 2261 37657 2295
rect 37657 2261 37691 2295
rect 37691 2261 37700 2295
rect 37648 2252 37700 2261
rect 10472 2150 10524 2202
rect 10536 2150 10588 2202
rect 10600 2150 10652 2202
rect 10664 2150 10716 2202
rect 10728 2150 10780 2202
rect 19994 2150 20046 2202
rect 20058 2150 20110 2202
rect 20122 2150 20174 2202
rect 20186 2150 20238 2202
rect 20250 2150 20302 2202
rect 29516 2150 29568 2202
rect 29580 2150 29632 2202
rect 29644 2150 29696 2202
rect 29708 2150 29760 2202
rect 29772 2150 29824 2202
rect 39038 2150 39090 2202
rect 39102 2150 39154 2202
rect 39166 2150 39218 2202
rect 39230 2150 39282 2202
rect 39294 2150 39346 2202
rect 3240 2048 3292 2100
rect 13820 2048 13872 2100
rect 23204 2048 23256 2100
rect 4712 1980 4764 2032
rect 7012 1980 7064 2032
rect 12348 1980 12400 2032
rect 29736 1980 29788 2032
rect 29920 2048 29972 2100
rect 35992 2048 36044 2100
rect 32588 1980 32640 2032
rect 5448 1912 5500 1964
rect 12164 1912 12216 1964
rect 16488 1912 16540 1964
rect 37556 1912 37608 1964
rect 6092 1844 6144 1896
rect 9496 1844 9548 1896
rect 13544 1844 13596 1896
rect 29644 1844 29696 1896
rect 29736 1844 29788 1896
rect 33508 1844 33560 1896
rect 6552 1776 6604 1828
rect 16764 1776 16816 1828
rect 24584 1776 24636 1828
rect 31668 1776 31720 1828
rect 12164 1708 12216 1760
rect 30380 1708 30432 1760
rect 14556 1640 14608 1692
rect 25504 1640 25556 1692
rect 29644 1640 29696 1692
rect 33600 1640 33652 1692
rect 4068 1572 4120 1624
rect 20720 1572 20772 1624
rect 8484 1504 8536 1556
rect 16212 1504 16264 1556
rect 2320 1300 2372 1352
rect 37372 1300 37424 1352
rect 7380 1232 7432 1284
rect 38568 1232 38620 1284
rect 6276 1164 6328 1216
rect 35164 1164 35216 1216
rect 11796 1096 11848 1148
rect 28908 1096 28960 1148
rect 1860 960 1912 1012
rect 3240 960 3292 1012
rect 2964 892 3016 944
rect 5172 892 5224 944
rect 11152 892 11204 944
rect 15476 892 15528 944
rect 15936 892 15988 944
rect 17408 892 17460 944
rect 21088 892 21140 944
rect 22560 892 22612 944
rect 29644 892 29696 944
rect 30748 892 30800 944
rect 31576 892 31628 944
rect 33140 892 33192 944
rect 33508 892 33560 944
rect 36636 892 36688 944
rect 36728 892 36780 944
rect 37648 892 37700 944
rect 5540 76 5592 128
rect 10232 76 10284 128
<< metal2 >>
rect 662 28354 718 29154
rect 1950 28506 2006 29154
rect 3882 28506 3938 29154
rect 1950 28478 2084 28506
rect 1950 28354 2006 28478
rect 676 26586 704 28354
rect 1030 27976 1086 27985
rect 1030 27911 1086 27920
rect 664 26580 716 26586
rect 664 26522 716 26528
rect 940 26036 992 26042
rect 940 25978 992 25984
rect 952 25945 980 25978
rect 938 25936 994 25945
rect 938 25871 994 25880
rect 1044 25498 1072 27911
rect 2056 26382 2084 28478
rect 3882 28478 4016 28506
rect 3882 28354 3938 28478
rect 2320 26852 2372 26858
rect 2320 26794 2372 26800
rect 2332 26450 2360 26794
rect 2320 26444 2372 26450
rect 2320 26386 2372 26392
rect 3988 26382 4016 28478
rect 5814 28354 5870 29154
rect 7746 28506 7802 29154
rect 9034 28506 9090 29154
rect 10966 28506 11022 29154
rect 12898 28506 12954 29154
rect 14830 28506 14886 29154
rect 7746 28478 8064 28506
rect 7746 28354 7802 28478
rect 5828 27146 5856 28354
rect 5828 27118 6132 27146
rect 5711 26684 6019 26693
rect 5711 26682 5717 26684
rect 5773 26682 5797 26684
rect 5853 26682 5877 26684
rect 5933 26682 5957 26684
rect 6013 26682 6019 26684
rect 5773 26630 5775 26682
rect 5955 26630 5957 26682
rect 5711 26628 5717 26630
rect 5773 26628 5797 26630
rect 5853 26628 5877 26630
rect 5933 26628 5957 26630
rect 6013 26628 6019 26630
rect 5711 26619 6019 26628
rect 6104 26382 6132 27118
rect 8036 26586 8064 28478
rect 9034 28478 9168 28506
rect 9034 28354 9090 28478
rect 8024 26580 8076 26586
rect 8024 26522 8076 26528
rect 9140 26382 9168 28478
rect 10966 28478 11376 28506
rect 10966 28354 11022 28478
rect 11348 26382 11376 28478
rect 12898 28478 13032 28506
rect 12898 28354 12954 28478
rect 13004 26382 13032 28478
rect 14830 28478 14964 28506
rect 14830 28354 14886 28478
rect 13084 26444 13136 26450
rect 13084 26386 13136 26392
rect 2044 26376 2096 26382
rect 3976 26376 4028 26382
rect 2044 26318 2096 26324
rect 3054 26344 3110 26353
rect 3976 26318 4028 26324
rect 6092 26376 6144 26382
rect 9128 26376 9180 26382
rect 6092 26318 6144 26324
rect 7930 26344 7986 26353
rect 3054 26279 3056 26288
rect 3108 26279 3110 26288
rect 9128 26318 9180 26324
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 7930 26279 7932 26288
rect 3056 26250 3108 26256
rect 7984 26279 7986 26288
rect 9404 26308 9456 26314
rect 7932 26250 7984 26256
rect 9404 26250 9456 26256
rect 2136 25900 2188 25906
rect 2136 25842 2188 25848
rect 1032 25492 1084 25498
rect 1032 25434 1084 25440
rect 940 24200 992 24206
rect 940 24142 992 24148
rect 952 23905 980 24142
rect 938 23896 994 23905
rect 938 23831 994 23840
rect 938 22536 994 22545
rect 938 22471 994 22480
rect 952 22438 980 22471
rect 940 22432 992 22438
rect 940 22374 992 22380
rect 940 20936 992 20942
rect 940 20878 992 20884
rect 952 20505 980 20878
rect 938 20496 994 20505
rect 938 20431 994 20440
rect 940 18624 992 18630
rect 940 18566 992 18572
rect 952 18465 980 18566
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 940 16516 992 16522
rect 940 16458 992 16464
rect 952 16425 980 16458
rect 938 16416 994 16425
rect 938 16351 994 16360
rect 1596 16114 1624 17138
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 940 15496 992 15502
rect 940 15438 992 15444
rect 952 15065 980 15438
rect 938 15056 994 15065
rect 938 14991 994 15000
rect 1596 13326 1624 16050
rect 1780 14618 1808 17682
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1676 14340 1728 14346
rect 1676 14282 1728 14288
rect 1688 13841 1716 14282
rect 1674 13832 1730 13841
rect 1674 13767 1730 13776
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 940 13184 992 13190
rect 940 13126 992 13132
rect 952 13025 980 13126
rect 938 13016 994 13025
rect 938 12951 994 12960
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1780 11762 1808 12378
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1872 11642 1900 16934
rect 2056 16590 2084 17614
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2042 15600 2098 15609
rect 2042 15535 2098 15544
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14414 1992 14758
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 2056 14006 2084 15535
rect 2148 14618 2176 25842
rect 8392 25832 8444 25838
rect 8392 25774 8444 25780
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 5711 25596 6019 25605
rect 5711 25594 5717 25596
rect 5773 25594 5797 25596
rect 5853 25594 5877 25596
rect 5933 25594 5957 25596
rect 6013 25594 6019 25596
rect 5773 25542 5775 25594
rect 5955 25542 5957 25594
rect 5711 25540 5717 25542
rect 5773 25540 5797 25542
rect 5853 25540 5877 25542
rect 5933 25540 5957 25542
rect 6013 25540 6019 25542
rect 5711 25531 6019 25540
rect 8300 25492 8352 25498
rect 8300 25434 8352 25440
rect 7932 25288 7984 25294
rect 7932 25230 7984 25236
rect 6184 25152 6236 25158
rect 6184 25094 6236 25100
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 5711 24508 6019 24517
rect 5711 24506 5717 24508
rect 5773 24506 5797 24508
rect 5853 24506 5877 24508
rect 5933 24506 5957 24508
rect 6013 24506 6019 24508
rect 5773 24454 5775 24506
rect 5955 24454 5957 24506
rect 5711 24452 5717 24454
rect 5773 24452 5797 24454
rect 5853 24452 5877 24454
rect 5933 24452 5957 24454
rect 6013 24452 6019 24454
rect 5711 24443 6019 24452
rect 6196 24274 6224 25094
rect 6184 24268 6236 24274
rect 6184 24210 6236 24216
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 2228 24132 2280 24138
rect 2228 24074 2280 24080
rect 6092 24132 6144 24138
rect 6092 24074 6144 24080
rect 2240 23594 2268 24074
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 2228 23588 2280 23594
rect 2228 23530 2280 23536
rect 2964 23520 3016 23526
rect 2964 23462 3016 23468
rect 2228 23248 2280 23254
rect 2228 23190 2280 23196
rect 2240 22778 2268 23190
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2240 19174 2268 20334
rect 2688 19848 2740 19854
rect 2688 19790 2740 19796
rect 2700 19378 2728 19790
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2228 19168 2280 19174
rect 2228 19110 2280 19116
rect 2240 18222 2268 19110
rect 2872 18692 2924 18698
rect 2872 18634 2924 18640
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2240 17134 2268 18158
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2780 17536 2832 17542
rect 2780 17478 2832 17484
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2240 16046 2268 17070
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2240 14890 2268 15982
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2332 14482 2360 14894
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2044 14000 2096 14006
rect 2044 13942 2096 13948
rect 2136 13864 2188 13870
rect 2188 13812 2268 13818
rect 2136 13806 2268 13812
rect 2148 13790 2268 13806
rect 2136 13456 2188 13462
rect 2136 13398 2188 13404
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2056 12850 2084 13262
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 1780 11614 1900 11642
rect 1780 11098 1808 11614
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11257 1900 11494
rect 1858 11248 1914 11257
rect 1858 11183 1914 11192
rect 940 11076 992 11082
rect 1780 11070 1900 11098
rect 940 11018 992 11024
rect 952 10985 980 11018
rect 938 10976 994 10985
rect 938 10911 994 10920
rect 1768 10056 1820 10062
rect 1688 10004 1768 10010
rect 1688 9998 1820 10004
rect 1688 9982 1808 9998
rect 1032 9920 1084 9926
rect 1032 9862 1084 9868
rect 20 8968 72 8974
rect 20 8910 72 8916
rect 938 8936 994 8945
rect 32 800 60 8910
rect 938 8871 994 8880
rect 952 8498 980 8871
rect 940 8492 992 8498
rect 940 8434 992 8440
rect 938 7576 994 7585
rect 938 7511 994 7520
rect 952 6322 980 7511
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 1044 5545 1072 9862
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1030 5536 1086 5545
rect 1030 5471 1086 5480
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 3505 980 5170
rect 1308 3528 1360 3534
rect 938 3496 994 3505
rect 1308 3470 1360 3476
rect 938 3431 994 3440
rect 1320 800 1348 3470
rect 1412 1465 1440 9522
rect 1688 7410 1716 9982
rect 1766 9480 1822 9489
rect 1766 9415 1822 9424
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1584 6180 1636 6186
rect 1584 6122 1636 6128
rect 1596 5710 1624 6122
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 5098 1624 5646
rect 1584 5092 1636 5098
rect 1584 5034 1636 5040
rect 1596 4622 1624 5034
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1596 4078 1624 4558
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1596 3058 1624 4014
rect 1688 3670 1716 7346
rect 1780 5370 1808 9415
rect 1872 6866 1900 11070
rect 1964 10742 1992 12650
rect 2056 12306 2084 12786
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 7818 1992 8366
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1872 4690 1900 6054
rect 1964 5914 1992 6666
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2056 5302 2084 11494
rect 2148 9042 2176 13398
rect 2240 12782 2268 13790
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2240 11898 2268 12718
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2424 10742 2452 17478
rect 2792 16697 2820 17478
rect 2778 16688 2834 16697
rect 2778 16623 2834 16632
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2700 16250 2728 16390
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2516 15706 2544 15982
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2700 15201 2728 15370
rect 2686 15192 2742 15201
rect 2686 15127 2742 15136
rect 2596 15088 2648 15094
rect 2596 15030 2648 15036
rect 2608 14618 2636 15030
rect 2700 14804 2728 15127
rect 2700 14776 2820 14804
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2226 10024 2282 10033
rect 2226 9959 2228 9968
rect 2280 9959 2282 9968
rect 2228 9930 2280 9936
rect 2332 9178 2360 10542
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2424 9110 2452 9454
rect 2412 9104 2464 9110
rect 2412 9046 2464 9052
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 2148 6730 2176 7754
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7478 2452 7686
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1780 2774 1808 3878
rect 1858 3632 1914 3641
rect 1858 3567 1860 3576
rect 1912 3567 1914 3576
rect 1860 3538 1912 3544
rect 1858 3224 1914 3233
rect 1858 3159 1914 3168
rect 1872 3126 1900 3159
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 2240 2774 2268 7142
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 5778 2360 6598
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2424 5030 2452 6666
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2516 4554 2544 13126
rect 2596 12232 2648 12238
rect 2792 12209 2820 14776
rect 2596 12174 2648 12180
rect 2778 12200 2834 12209
rect 2608 10130 2636 12174
rect 2778 12135 2834 12144
rect 2688 12096 2740 12102
rect 2884 12050 2912 18634
rect 2976 18358 3004 23462
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 3068 21078 3096 21830
rect 3056 21072 3108 21078
rect 3056 21014 3108 21020
rect 2964 18352 3016 18358
rect 2964 18294 3016 18300
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2688 12038 2740 12044
rect 2700 11558 2728 12038
rect 2792 12022 2912 12050
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2792 10554 2820 12022
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2884 11150 2912 11834
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2884 10674 2912 11086
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2792 10526 2912 10554
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2608 9761 2636 9930
rect 2594 9752 2650 9761
rect 2594 9687 2650 9696
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2608 6730 2636 8978
rect 2700 7818 2728 10202
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2792 7993 2820 8434
rect 2778 7984 2834 7993
rect 2778 7919 2834 7928
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2792 7274 2820 7822
rect 2780 7268 2832 7274
rect 2780 7210 2832 7216
rect 2778 7168 2834 7177
rect 2778 7103 2834 7112
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2700 5681 2728 6190
rect 2686 5672 2742 5681
rect 2686 5607 2742 5616
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2608 3738 2636 5102
rect 2792 4321 2820 7103
rect 2884 6882 2912 10526
rect 2976 9178 3004 15846
rect 3068 15450 3096 21014
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3160 15994 3188 16526
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 3252 16182 3280 16390
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 3160 15966 3280 15994
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3160 15570 3188 15846
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 3068 15422 3188 15450
rect 3056 15360 3108 15366
rect 3054 15328 3056 15337
rect 3108 15328 3110 15337
rect 3054 15263 3110 15272
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 3068 14482 3096 14758
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3160 14346 3188 15422
rect 3252 15042 3280 15966
rect 3344 15570 3372 22034
rect 3422 17640 3478 17649
rect 3422 17575 3478 17584
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3252 15014 3372 15042
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3344 13410 3372 15014
rect 3436 14006 3464 17575
rect 3424 14000 3476 14006
rect 3424 13942 3476 13948
rect 3344 13382 3464 13410
rect 3332 13320 3384 13326
rect 3330 13288 3332 13297
rect 3384 13288 3386 13297
rect 3330 13223 3386 13232
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2976 7002 3004 8026
rect 3068 7410 3096 11222
rect 3160 11218 3188 12242
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3160 8498 3188 8978
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3160 7410 3188 7822
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 3054 6896 3110 6905
rect 2884 6854 3004 6882
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2884 6254 2912 6666
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2778 4312 2834 4321
rect 2778 4247 2834 4256
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2792 3534 2820 4247
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 3466 2912 6190
rect 2976 4214 3004 6854
rect 3054 6831 3110 6840
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 3068 4078 3096 6831
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6497 3188 6598
rect 3146 6488 3202 6497
rect 3146 6423 3202 6432
rect 3252 5642 3280 12038
rect 3436 11898 3464 13382
rect 3528 12918 3556 22918
rect 3700 22432 3752 22438
rect 3700 22374 3752 22380
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3620 15706 3648 21830
rect 3712 18358 3740 22374
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3620 14346 3648 15642
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3712 13870 3740 14350
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3620 12442 3648 12650
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3514 12200 3570 12209
rect 3514 12135 3570 12144
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3344 8294 3372 8570
rect 3436 8537 3464 11154
rect 3422 8528 3478 8537
rect 3422 8463 3478 8472
rect 3436 8430 3464 8463
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3332 8288 3384 8294
rect 3384 8248 3464 8276
rect 3332 8230 3384 8236
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3344 7546 3372 8026
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3436 6458 3464 8248
rect 3528 6497 3556 12135
rect 3712 9042 3740 13398
rect 3804 12918 3832 23122
rect 4068 23112 4120 23118
rect 4172 23066 4200 23666
rect 4896 23656 4948 23662
rect 4896 23598 4948 23604
rect 4120 23060 4200 23066
rect 4068 23054 4200 23060
rect 4080 23038 4200 23054
rect 4068 22636 4120 22642
rect 4172 22624 4200 23038
rect 4712 23044 4764 23050
rect 4712 22986 4764 22992
rect 4120 22596 4200 22624
rect 4068 22578 4120 22584
rect 3976 22500 4028 22506
rect 3976 22442 4028 22448
rect 3988 22166 4016 22442
rect 3976 22160 4028 22166
rect 3976 22102 4028 22108
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 3896 20398 3924 21830
rect 4080 21690 4108 22578
rect 4252 21956 4304 21962
rect 4252 21898 4304 21904
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4080 20942 4108 21626
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 3884 19440 3936 19446
rect 3884 19382 3936 19388
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3896 12434 3924 19382
rect 3988 17202 4016 20742
rect 4172 20262 4200 21830
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4172 19990 4200 20198
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 4264 19836 4292 21898
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4448 21690 4476 21830
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 4172 19808 4292 19836
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3988 14958 4016 15438
rect 4172 15434 4200 19808
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 4264 15094 4292 19654
rect 4448 18766 4476 19654
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4356 16454 4384 17070
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4448 16454 4476 16934
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4540 16114 4568 21490
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4632 15994 4660 16594
rect 4448 15966 4660 15994
rect 4342 15464 4398 15473
rect 4342 15399 4398 15408
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3988 14482 4016 14894
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 4356 14414 4384 15399
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3804 12406 3924 12434
rect 3804 11762 3832 12406
rect 3988 12238 4016 13874
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13530 4108 13670
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4448 13190 4476 15966
rect 4526 15872 4582 15881
rect 4526 15807 4582 15816
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4448 12918 4476 13126
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4540 12782 4568 15807
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4632 13920 4660 15506
rect 4724 15434 4752 22986
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 4816 22234 4844 22374
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 4908 22166 4936 23598
rect 5711 23420 6019 23429
rect 5711 23418 5717 23420
rect 5773 23418 5797 23420
rect 5853 23418 5877 23420
rect 5933 23418 5957 23420
rect 6013 23418 6019 23420
rect 5773 23366 5775 23418
rect 5955 23366 5957 23418
rect 5711 23364 5717 23366
rect 5773 23364 5797 23366
rect 5853 23364 5877 23366
rect 5933 23364 5957 23366
rect 6013 23364 6019 23366
rect 5711 23355 6019 23364
rect 5632 22432 5684 22438
rect 5632 22374 5684 22380
rect 4896 22160 4948 22166
rect 4896 22102 4948 22108
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4816 15337 4844 16934
rect 4908 16658 4936 22102
rect 5540 20868 5592 20874
rect 5540 20810 5592 20816
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 5184 17202 5212 19178
rect 5552 17218 5580 20810
rect 5644 19922 5672 22374
rect 5711 22332 6019 22341
rect 5711 22330 5717 22332
rect 5773 22330 5797 22332
rect 5853 22330 5877 22332
rect 5933 22330 5957 22332
rect 6013 22330 6019 22332
rect 5773 22278 5775 22330
rect 5955 22278 5957 22330
rect 5711 22276 5717 22278
rect 5773 22276 5797 22278
rect 5853 22276 5877 22278
rect 5933 22276 5957 22278
rect 6013 22276 6019 22278
rect 5711 22267 6019 22276
rect 5711 21244 6019 21253
rect 5711 21242 5717 21244
rect 5773 21242 5797 21244
rect 5853 21242 5877 21244
rect 5933 21242 5957 21244
rect 6013 21242 6019 21244
rect 5773 21190 5775 21242
rect 5955 21190 5957 21242
rect 5711 21188 5717 21190
rect 5773 21188 5797 21190
rect 5853 21188 5877 21190
rect 5933 21188 5957 21190
rect 6013 21188 6019 21190
rect 5711 21179 6019 21188
rect 5711 20156 6019 20165
rect 5711 20154 5717 20156
rect 5773 20154 5797 20156
rect 5853 20154 5877 20156
rect 5933 20154 5957 20156
rect 6013 20154 6019 20156
rect 5773 20102 5775 20154
rect 5955 20102 5957 20154
rect 5711 20100 5717 20102
rect 5773 20100 5797 20102
rect 5853 20100 5877 20102
rect 5933 20100 5957 20102
rect 6013 20100 6019 20102
rect 5711 20091 6019 20100
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5644 18766 5672 19246
rect 6012 19242 6040 19994
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 6104 19174 6132 24074
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 6196 19854 6224 22374
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 5711 19068 6019 19077
rect 5711 19066 5717 19068
rect 5773 19066 5797 19068
rect 5853 19066 5877 19068
rect 5933 19066 5957 19068
rect 6013 19066 6019 19068
rect 5773 19014 5775 19066
rect 5955 19014 5957 19066
rect 5711 19012 5717 19014
rect 5773 19012 5797 19014
rect 5853 19012 5877 19014
rect 5933 19012 5957 19014
rect 6013 19012 6019 19014
rect 5711 19003 6019 19012
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5460 17190 5580 17218
rect 5184 17105 5212 17138
rect 5170 17096 5226 17105
rect 5080 17060 5132 17066
rect 5354 17096 5410 17105
rect 5170 17031 5226 17040
rect 5276 17054 5354 17082
rect 5080 17002 5132 17008
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4802 15328 4858 15337
rect 4802 15263 4858 15272
rect 5000 15162 5028 16390
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 4908 15065 4936 15098
rect 4894 15056 4950 15065
rect 4894 14991 4950 15000
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5000 14521 5028 14554
rect 4986 14512 5042 14521
rect 4986 14447 5042 14456
rect 4632 13892 5028 13920
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3896 11354 3924 12106
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3988 11150 4016 12174
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4264 11082 4292 11494
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 3896 10962 3924 11018
rect 3896 10934 4016 10962
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3804 8974 3832 10406
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3606 7712 3662 7721
rect 3606 7647 3662 7656
rect 3620 7478 3648 7647
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3514 6488 3570 6497
rect 3424 6452 3476 6458
rect 3514 6423 3570 6432
rect 3424 6394 3476 6400
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3344 4690 3372 6326
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3436 4162 3464 6122
rect 3620 4434 3648 7278
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3712 5778 3740 6190
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3698 5672 3754 5681
rect 3698 5607 3754 5616
rect 3712 4622 3740 5607
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3620 4406 3740 4434
rect 3344 4134 3464 4162
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 3344 2774 3372 4134
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3436 3126 3464 4014
rect 3514 3632 3570 3641
rect 3514 3567 3516 3576
rect 3568 3567 3570 3576
rect 3516 3538 3568 3544
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3712 2990 3740 4406
rect 3804 3058 3832 8910
rect 3896 8022 3924 10542
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 5098 3924 7686
rect 3988 7562 4016 10934
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4172 9518 4200 9862
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4068 9172 4120 9178
rect 4264 9160 4292 9454
rect 4068 9114 4120 9120
rect 4172 9132 4292 9160
rect 4080 8673 4108 9114
rect 4066 8664 4122 8673
rect 4066 8599 4122 8608
rect 4066 7576 4122 7585
rect 3988 7534 4066 7562
rect 4066 7511 4122 7520
rect 4080 6662 4108 7511
rect 4172 6730 4200 9132
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4264 8634 4292 8978
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4264 8498 4292 8570
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4356 7886 4384 11290
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4448 8090 4476 9930
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4540 9382 4568 9862
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4632 8922 4660 13126
rect 4894 11656 4950 11665
rect 4894 11591 4950 11600
rect 4908 10130 4936 11591
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4540 8894 4660 8922
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4448 7410 4476 7482
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4342 7304 4398 7313
rect 4342 7239 4398 7248
rect 4356 6866 4384 7239
rect 4448 6934 4476 7346
rect 4436 6928 4488 6934
rect 4540 6905 4568 8894
rect 4618 8664 4674 8673
rect 4618 8599 4674 8608
rect 4632 8566 4660 8599
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4436 6870 4488 6876
rect 4526 6896 4582 6905
rect 4344 6860 4396 6866
rect 4526 6831 4582 6840
rect 4344 6802 4396 6808
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3988 6390 4016 6598
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 4080 6254 4108 6598
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4172 5658 4200 6666
rect 4264 6458 4292 6666
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 3988 5630 4200 5658
rect 3988 5574 4016 5630
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3974 4040 4030 4049
rect 3974 3975 4030 3984
rect 3988 3738 4016 3975
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 1780 2746 1900 2774
rect 2240 2746 2360 2774
rect 3344 2746 3648 2774
rect 1398 1456 1454 1465
rect 1398 1391 1454 1400
rect 1872 1018 1900 2746
rect 2332 1358 2360 2746
rect 3620 2514 3648 2746
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2320 1352 2372 1358
rect 2320 1294 2372 1300
rect 1860 1012 1912 1018
rect 1860 954 1912 960
rect 2976 950 3004 2382
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 3252 2106 3280 2314
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 4080 1630 4108 5510
rect 4264 4622 4292 6394
rect 4356 6236 4384 6802
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4448 6390 4476 6734
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4356 6208 4476 6236
rect 4342 5808 4398 5817
rect 4342 5743 4398 5752
rect 4356 5302 4384 5743
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4172 3126 4200 4558
rect 4356 4162 4384 5238
rect 4264 4134 4384 4162
rect 4264 3534 4292 4134
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4172 2378 4200 3062
rect 4356 3058 4384 3946
rect 4448 3602 4476 6208
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5710 4568 6054
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4526 5536 4582 5545
rect 4526 5471 4582 5480
rect 4540 4826 4568 5471
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4632 4486 4660 7890
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4526 4176 4582 4185
rect 4526 4111 4582 4120
rect 4540 4078 4568 4111
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4632 3534 4660 4422
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4724 2650 4752 7754
rect 4816 7546 4844 8978
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4802 7440 4858 7449
rect 4802 7375 4804 7384
rect 4856 7375 4858 7384
rect 4804 7346 4856 7352
rect 4908 7313 4936 10066
rect 5000 8906 5028 13892
rect 5092 11665 5120 17002
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5184 14346 5212 15982
rect 5276 14890 5304 17054
rect 5354 17031 5410 17040
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5368 16794 5396 16934
rect 5460 16794 5488 17190
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 5368 13818 5396 14826
rect 5460 13938 5488 16390
rect 5552 15094 5580 17070
rect 5644 16590 5672 18702
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5736 18426 5764 18566
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5711 17980 6019 17989
rect 5711 17978 5717 17980
rect 5773 17978 5797 17980
rect 5853 17978 5877 17980
rect 5933 17978 5957 17980
rect 6013 17978 6019 17980
rect 5773 17926 5775 17978
rect 5955 17926 5957 17978
rect 5711 17924 5717 17926
rect 5773 17924 5797 17926
rect 5853 17924 5877 17926
rect 5933 17924 5957 17926
rect 6013 17924 6019 17926
rect 5711 17915 6019 17924
rect 5711 16892 6019 16901
rect 5711 16890 5717 16892
rect 5773 16890 5797 16892
rect 5853 16890 5877 16892
rect 5933 16890 5957 16892
rect 6013 16890 6019 16892
rect 5773 16838 5775 16890
rect 5955 16838 5957 16890
rect 5711 16836 5717 16838
rect 5773 16836 5797 16838
rect 5853 16836 5877 16838
rect 5933 16836 5957 16838
rect 6013 16836 6019 16838
rect 5711 16827 6019 16836
rect 6288 16810 6316 22918
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 6196 16782 6316 16810
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5644 16182 5672 16526
rect 6012 16402 6040 16730
rect 6012 16374 6132 16402
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 5644 15502 5672 16118
rect 5711 15804 6019 15813
rect 5711 15802 5717 15804
rect 5773 15802 5797 15804
rect 5853 15802 5877 15804
rect 5933 15802 5957 15804
rect 6013 15802 6019 15804
rect 5773 15750 5775 15802
rect 5955 15750 5957 15802
rect 5711 15748 5717 15750
rect 5773 15748 5797 15750
rect 5853 15748 5877 15750
rect 5933 15748 5957 15750
rect 6013 15748 6019 15750
rect 5711 15739 6019 15748
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5632 15088 5684 15094
rect 5632 15030 5684 15036
rect 5552 14822 5580 15030
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5540 13864 5592 13870
rect 5368 13812 5540 13818
rect 5368 13806 5592 13812
rect 5368 13790 5580 13806
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5184 12850 5212 13262
rect 5368 13258 5396 13790
rect 5644 13734 5672 15030
rect 5711 14716 6019 14725
rect 5711 14714 5717 14716
rect 5773 14714 5797 14716
rect 5853 14714 5877 14716
rect 5933 14714 5957 14716
rect 6013 14714 6019 14716
rect 5773 14662 5775 14714
rect 5955 14662 5957 14714
rect 5711 14660 5717 14662
rect 5773 14660 5797 14662
rect 5853 14660 5877 14662
rect 5933 14660 5957 14662
rect 6013 14660 6019 14662
rect 5711 14651 6019 14660
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5711 13628 6019 13637
rect 5711 13626 5717 13628
rect 5773 13626 5797 13628
rect 5853 13626 5877 13628
rect 5933 13626 5957 13628
rect 6013 13626 6019 13628
rect 5773 13574 5775 13626
rect 5955 13574 5957 13626
rect 5711 13572 5717 13574
rect 5773 13572 5797 13574
rect 5853 13572 5877 13574
rect 5933 13572 5957 13574
rect 6013 13572 6019 13574
rect 5711 13563 6019 13572
rect 6104 13512 6132 16374
rect 6012 13484 6132 13512
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5264 12640 5316 12646
rect 5262 12608 5264 12617
rect 5316 12608 5318 12617
rect 5262 12543 5318 12552
rect 5460 11898 5488 13330
rect 6012 13190 6040 13484
rect 6196 13410 6224 16782
rect 6380 15094 6408 20946
rect 6564 20466 6592 24210
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6656 23866 6684 24074
rect 7208 23866 7236 25094
rect 7668 24070 7696 25094
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6736 22976 6788 22982
rect 6736 22918 6788 22924
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6564 18766 6592 20402
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6656 15502 6684 17614
rect 6748 17218 6776 22918
rect 6840 17338 6868 23462
rect 6932 18329 6960 23666
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 7024 22506 7052 23122
rect 7668 22710 7696 24006
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 7656 22704 7708 22710
rect 7656 22646 7708 22652
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 6918 18320 6974 18329
rect 6918 18255 6974 18264
rect 6932 18222 6960 18255
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 6748 17190 6868 17218
rect 6840 16998 6868 17190
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6840 16182 6868 16934
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6656 15337 6684 15438
rect 6642 15328 6698 15337
rect 6642 15263 6698 15272
rect 6368 15088 6420 15094
rect 6368 15030 6420 15036
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6104 13382 6224 13410
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6104 12986 6132 13382
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 6196 12986 6224 13194
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12238 5672 12786
rect 5711 12540 6019 12549
rect 5711 12538 5717 12540
rect 5773 12538 5797 12540
rect 5853 12538 5877 12540
rect 5933 12538 5957 12540
rect 6013 12538 6019 12540
rect 5773 12486 5775 12538
rect 5955 12486 5957 12538
rect 5711 12484 5717 12486
rect 5773 12484 5797 12486
rect 5853 12484 5877 12486
rect 5933 12484 5957 12486
rect 6013 12484 6019 12486
rect 5711 12475 6019 12484
rect 6288 12434 6316 14758
rect 6748 14618 6776 14962
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 7102 14512 7158 14521
rect 7012 14476 7064 14482
rect 7102 14447 7158 14456
rect 7012 14418 7064 14424
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6564 14074 6592 14282
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6656 14074 6684 14214
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6564 13394 6592 14010
rect 6748 13977 6776 14214
rect 6734 13968 6790 13977
rect 6734 13903 6790 13912
rect 6644 13728 6696 13734
rect 6642 13696 6644 13705
rect 6696 13696 6698 13705
rect 6642 13631 6698 13640
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6104 12406 6316 12434
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5078 11656 5134 11665
rect 5078 11591 5134 11600
rect 5368 11286 5396 11834
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 5080 8832 5132 8838
rect 5000 8780 5080 8786
rect 5000 8774 5132 8780
rect 5000 8758 5120 8774
rect 4894 7304 4950 7313
rect 4894 7239 4950 7248
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4816 3641 4844 6802
rect 4896 5636 4948 5642
rect 4896 5578 4948 5584
rect 4908 4826 4936 5578
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5000 4298 5028 8758
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5092 7206 5120 7686
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5184 6361 5212 9998
rect 5276 7324 5304 10746
rect 5368 10266 5396 10746
rect 5446 10568 5502 10577
rect 5446 10503 5502 10512
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5460 9586 5488 10503
rect 5552 10146 5580 11630
rect 5644 11218 5672 11698
rect 5828 11694 5856 12242
rect 5816 11688 5868 11694
rect 5814 11656 5816 11665
rect 5868 11656 5870 11665
rect 5814 11591 5870 11600
rect 5711 11452 6019 11461
rect 5711 11450 5717 11452
rect 5773 11450 5797 11452
rect 5853 11450 5877 11452
rect 5933 11450 5957 11452
rect 6013 11450 6019 11452
rect 5773 11398 5775 11450
rect 5955 11398 5957 11450
rect 5711 11396 5717 11398
rect 5773 11396 5797 11398
rect 5853 11396 5877 11398
rect 5933 11396 5957 11398
rect 6013 11396 6019 11398
rect 5711 11387 6019 11396
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5644 10266 5672 11018
rect 5724 10736 5776 10742
rect 5722 10704 5724 10713
rect 5776 10704 5778 10713
rect 5722 10639 5778 10648
rect 6012 10538 6040 11222
rect 6104 11014 6132 12406
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 5711 10364 6019 10373
rect 5711 10362 5717 10364
rect 5773 10362 5797 10364
rect 5853 10362 5877 10364
rect 5933 10362 5957 10364
rect 6013 10362 6019 10364
rect 5773 10310 5775 10362
rect 5955 10310 5957 10362
rect 5711 10308 5717 10310
rect 5773 10308 5797 10310
rect 5853 10308 5877 10310
rect 5933 10308 5957 10310
rect 6013 10308 6019 10310
rect 5711 10299 6019 10308
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5552 10118 5672 10146
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5552 9654 5580 9998
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5446 8528 5502 8537
rect 5446 8463 5502 8472
rect 5276 7296 5396 7324
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5170 6352 5226 6361
rect 5170 6287 5226 6296
rect 5276 5914 5304 7142
rect 5368 6633 5396 7296
rect 5354 6624 5410 6633
rect 5354 6559 5410 6568
rect 5460 6236 5488 8463
rect 5552 6662 5580 9318
rect 5644 8974 5672 10118
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5828 9586 5856 10066
rect 6104 9994 6132 10950
rect 6092 9988 6144 9994
rect 6092 9930 6144 9936
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 5711 9276 6019 9285
rect 5711 9274 5717 9276
rect 5773 9274 5797 9276
rect 5853 9274 5877 9276
rect 5933 9274 5957 9276
rect 6013 9274 6019 9276
rect 5773 9222 5775 9274
rect 5955 9222 5957 9274
rect 5711 9220 5717 9222
rect 5773 9220 5797 9222
rect 5853 9220 5877 9222
rect 5933 9220 5957 9222
rect 6013 9220 6019 9222
rect 5711 9211 6019 9220
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5644 8294 5672 8910
rect 5632 8288 5684 8294
rect 6012 8276 6040 9114
rect 6104 9110 6132 9318
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6012 8248 6132 8276
rect 5632 8230 5684 8236
rect 5644 7886 5672 8230
rect 5711 8188 6019 8197
rect 5711 8186 5717 8188
rect 5773 8186 5797 8188
rect 5853 8186 5877 8188
rect 5933 8186 5957 8188
rect 6013 8186 6019 8188
rect 5773 8134 5775 8186
rect 5955 8134 5957 8186
rect 5711 8132 5717 8134
rect 5773 8132 5797 8134
rect 5853 8132 5877 8134
rect 5933 8132 5957 8134
rect 6013 8132 6019 8134
rect 5711 8123 6019 8132
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5644 7206 5672 7822
rect 5722 7576 5778 7585
rect 5722 7511 5778 7520
rect 5736 7342 5764 7511
rect 5724 7336 5776 7342
rect 5816 7336 5868 7342
rect 5724 7278 5776 7284
rect 5814 7304 5816 7313
rect 5868 7304 5870 7313
rect 5814 7239 5870 7248
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5711 7100 6019 7109
rect 5711 7098 5717 7100
rect 5773 7098 5797 7100
rect 5853 7098 5877 7100
rect 5933 7098 5957 7100
rect 6013 7098 6019 7100
rect 5773 7046 5775 7098
rect 5955 7046 5957 7098
rect 5711 7044 5717 7046
rect 5773 7044 5797 7046
rect 5853 7044 5877 7046
rect 5933 7044 5957 7046
rect 6013 7044 6019 7046
rect 5711 7035 6019 7044
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5460 6208 5580 6236
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5092 4486 5120 4762
rect 5184 4690 5212 5510
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5184 4298 5212 4422
rect 5000 4270 5212 4298
rect 5184 4214 5212 4270
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 4802 3632 4858 3641
rect 4802 3567 4858 3576
rect 5184 3398 5212 4150
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5276 3194 5304 5170
rect 5354 5128 5410 5137
rect 5354 5063 5410 5072
rect 5368 3942 5396 5063
rect 5460 4282 5488 6054
rect 5552 4690 5580 6208
rect 5711 6012 6019 6021
rect 5711 6010 5717 6012
rect 5773 6010 5797 6012
rect 5853 6010 5877 6012
rect 5933 6010 5957 6012
rect 6013 6010 6019 6012
rect 5773 5958 5775 6010
rect 5955 5958 5957 6010
rect 5711 5956 5717 5958
rect 5773 5956 5797 5958
rect 5853 5956 5877 5958
rect 5933 5956 5957 5958
rect 6013 5956 6019 5958
rect 5711 5947 6019 5956
rect 5998 5400 6054 5409
rect 6104 5370 6132 8248
rect 6196 5642 6224 12038
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11286 6316 11494
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6380 11234 6408 13126
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6472 11830 6500 12038
rect 6656 11898 6684 13631
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6380 11206 6500 11234
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6288 10062 6316 11086
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6366 9752 6422 9761
rect 6366 9687 6422 9696
rect 6380 9654 6408 9687
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6288 8634 6316 9454
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6288 7954 6316 8570
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6202 6316 7142
rect 6380 6322 6408 8842
rect 6472 8401 6500 11206
rect 6748 10742 6776 13903
rect 7024 13870 7052 14418
rect 7116 14278 7144 14447
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7208 13734 7236 14350
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7288 13524 7340 13530
rect 7116 13484 7288 13512
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6840 11150 6868 11766
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6840 10588 6868 10950
rect 6932 10674 6960 13330
rect 7010 12608 7066 12617
rect 7010 12543 7066 12552
rect 7024 12306 7052 12543
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7010 11928 7066 11937
rect 7010 11863 7066 11872
rect 7024 11762 7052 11863
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6748 10560 6868 10588
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6458 8392 6514 8401
rect 6458 8327 6514 8336
rect 6460 7472 6512 7478
rect 6564 7460 6592 10066
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6512 7432 6592 7460
rect 6460 7414 6512 7420
rect 6564 7206 6592 7432
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6472 6866 6592 6882
rect 6460 6860 6592 6866
rect 6512 6854 6592 6860
rect 6460 6802 6512 6808
rect 6458 6760 6514 6769
rect 6458 6695 6460 6704
rect 6512 6695 6514 6704
rect 6460 6666 6512 6672
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6288 6174 6408 6202
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6288 5522 6316 5782
rect 6196 5494 6316 5522
rect 5998 5335 6054 5344
rect 6092 5364 6144 5370
rect 6012 5302 6040 5335
rect 6092 5306 6144 5312
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 5711 4924 6019 4933
rect 5711 4922 5717 4924
rect 5773 4922 5797 4924
rect 5853 4922 5877 4924
rect 5933 4922 5957 4924
rect 6013 4922 6019 4924
rect 5773 4870 5775 4922
rect 5955 4870 5957 4922
rect 5711 4868 5717 4870
rect 5773 4868 5797 4870
rect 5853 4868 5877 4870
rect 5933 4868 5957 4870
rect 6013 4868 6019 4870
rect 5711 4859 6019 4868
rect 6090 4856 6146 4865
rect 6090 4791 6146 4800
rect 6104 4758 6132 4791
rect 6092 4752 6144 4758
rect 5814 4720 5870 4729
rect 5540 4684 5592 4690
rect 6092 4694 6144 4700
rect 5814 4655 5870 4664
rect 5540 4626 5592 4632
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5644 3942 5672 4082
rect 5736 4049 5764 4490
rect 5828 4078 5856 4655
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5920 4214 5948 4558
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 5816 4072 5868 4078
rect 5722 4040 5778 4049
rect 5908 4072 5960 4078
rect 5816 4014 5868 4020
rect 5906 4040 5908 4049
rect 5960 4040 5962 4049
rect 5722 3975 5778 3984
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5632 3936 5684 3942
rect 5828 3924 5856 4014
rect 5906 3975 5962 3984
rect 5828 3896 6132 3924
rect 5632 3878 5684 3884
rect 5711 3836 6019 3845
rect 5711 3834 5717 3836
rect 5773 3834 5797 3836
rect 5853 3834 5877 3836
rect 5933 3834 5957 3836
rect 6013 3834 6019 3836
rect 5773 3782 5775 3834
rect 5955 3782 5957 3834
rect 5711 3780 5717 3782
rect 5773 3780 5797 3782
rect 5853 3780 5877 3782
rect 5933 3780 5957 3782
rect 6013 3780 6019 3782
rect 5711 3771 6019 3780
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4816 2961 4844 2994
rect 4802 2952 4858 2961
rect 4802 2887 4858 2896
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4816 2446 4844 2887
rect 5644 2514 5672 3538
rect 6012 3505 6040 3538
rect 5998 3496 6054 3505
rect 5998 3431 6054 3440
rect 5722 3360 5778 3369
rect 5722 3295 5778 3304
rect 5736 3194 5764 3295
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 6104 3126 6132 3896
rect 6092 3120 6144 3126
rect 5722 3088 5778 3097
rect 6092 3062 6144 3068
rect 5722 3023 5724 3032
rect 5776 3023 5778 3032
rect 5724 2994 5776 3000
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 5711 2748 6019 2757
rect 5711 2746 5717 2748
rect 5773 2746 5797 2748
rect 5853 2746 5877 2748
rect 5933 2746 5957 2748
rect 6013 2746 6019 2748
rect 5773 2694 5775 2746
rect 5955 2694 5957 2746
rect 5711 2692 5717 2694
rect 5773 2692 5797 2694
rect 5853 2692 5877 2694
rect 5933 2692 5957 2694
rect 6013 2692 6019 2694
rect 5711 2683 6019 2692
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 4724 2038 4752 2314
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 5460 1970 5488 2382
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5448 1964 5500 1970
rect 5448 1906 5500 1912
rect 4068 1624 4120 1630
rect 4068 1566 4120 1572
rect 3240 1012 3292 1018
rect 3240 954 3292 960
rect 2964 944 3016 950
rect 2964 886 3016 892
rect 3252 800 3280 954
rect 5172 944 5224 950
rect 5172 886 5224 892
rect 5184 800 5212 886
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 5170 0 5226 800
rect 5552 134 5580 2246
rect 6104 1902 6132 2926
rect 6196 2446 6224 5494
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 6092 1896 6144 1902
rect 6092 1838 6144 1844
rect 6288 1222 6316 3606
rect 6380 3398 6408 6174
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6472 2514 6500 6326
rect 6564 5710 6592 6854
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6564 5166 6592 5646
rect 6656 5642 6684 9862
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6564 4690 6592 5102
rect 6642 4856 6698 4865
rect 6642 4791 6698 4800
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6656 4264 6684 4791
rect 6564 4236 6684 4264
rect 6564 4078 6592 4236
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6564 1834 6592 3606
rect 6656 2961 6684 4082
rect 6748 3942 6776 10560
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6840 9518 6868 9998
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6840 8634 6868 8774
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6932 8514 6960 9862
rect 7024 8673 7052 11494
rect 7116 10470 7144 13484
rect 7288 13466 7340 13472
rect 7286 12880 7342 12889
rect 7286 12815 7342 12824
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7208 10112 7236 12650
rect 7300 11762 7328 12815
rect 7392 12753 7420 17274
rect 7760 17270 7788 23802
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7760 16046 7788 16526
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7470 13832 7526 13841
rect 7470 13767 7526 13776
rect 7484 13462 7512 13767
rect 7472 13456 7524 13462
rect 7472 13398 7524 13404
rect 7576 12850 7604 15438
rect 7852 14940 7880 23666
rect 7944 15162 7972 25230
rect 8312 24410 8340 25434
rect 8404 25362 8432 25774
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8484 24200 8536 24206
rect 8484 24142 8536 24148
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 8128 23186 8156 23666
rect 8208 23656 8260 23662
rect 8208 23598 8260 23604
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 8220 22574 8248 23598
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8206 17776 8262 17785
rect 8206 17711 8262 17720
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 8036 15042 8064 17138
rect 8220 15706 8248 17711
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8208 15360 8260 15366
rect 8300 15360 8352 15366
rect 8208 15302 8260 15308
rect 8298 15328 8300 15337
rect 8352 15328 8354 15337
rect 7760 14912 7880 14940
rect 7944 15014 8064 15042
rect 7760 13394 7788 14912
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7760 12986 7788 13330
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7472 12776 7524 12782
rect 7378 12744 7434 12753
rect 7472 12718 7524 12724
rect 7378 12679 7434 12688
rect 7378 12200 7434 12209
rect 7378 12135 7380 12144
rect 7432 12135 7434 12144
rect 7380 12106 7432 12112
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7392 11694 7420 12106
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7484 11234 7512 12718
rect 7576 12220 7604 12786
rect 7760 12617 7788 12922
rect 7852 12918 7880 13194
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7746 12608 7802 12617
rect 7746 12543 7802 12552
rect 7748 12232 7800 12238
rect 7576 12192 7748 12220
rect 7748 12174 7800 12180
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7852 11898 7880 12106
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7484 11206 7604 11234
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7378 10704 7434 10713
rect 7378 10639 7434 10648
rect 7208 10084 7328 10112
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7116 9722 7144 9930
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7208 9466 7236 9862
rect 7116 9438 7236 9466
rect 7116 9042 7144 9438
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7208 8838 7236 9318
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7010 8664 7066 8673
rect 7010 8599 7066 8608
rect 6840 8498 6960 8514
rect 6828 8492 6960 8498
rect 6880 8486 6960 8492
rect 7102 8528 7158 8537
rect 7102 8463 7158 8472
rect 6828 8434 6880 8440
rect 6840 8294 6868 8434
rect 7116 8430 7144 8463
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 7104 7948 7156 7954
rect 7208 7936 7236 8366
rect 7156 7908 7236 7936
rect 7104 7890 7156 7896
rect 7116 7410 7144 7890
rect 7300 7818 7328 10084
rect 7392 9674 7420 10639
rect 7484 9874 7512 11086
rect 7576 10554 7604 11206
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7668 10674 7696 11154
rect 7760 11150 7788 11562
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7576 10526 7696 10554
rect 7484 9846 7604 9874
rect 7392 9646 7512 9674
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7392 9178 7420 9454
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7484 8566 7512 9646
rect 7576 9382 7604 9846
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7576 8974 7604 9318
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7472 8560 7524 8566
rect 7668 8537 7696 10526
rect 7760 9178 7788 11086
rect 7852 9926 7880 11834
rect 7944 11762 7972 15014
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8022 13968 8078 13977
rect 8022 13903 8024 13912
rect 8076 13903 8078 13912
rect 8024 13874 8076 13880
rect 8024 13728 8076 13734
rect 8024 13670 8076 13676
rect 8036 13530 8064 13670
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12986 8064 13126
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8022 12744 8078 12753
rect 8022 12679 8078 12688
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8036 10742 8064 12679
rect 8128 11801 8156 14894
rect 8220 13977 8248 15302
rect 8298 15263 8354 15272
rect 8496 15201 8524 24142
rect 8944 24064 8996 24070
rect 8944 24006 8996 24012
rect 8956 23322 8984 24006
rect 8944 23316 8996 23322
rect 8944 23258 8996 23264
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8588 15858 8616 16186
rect 8666 16144 8722 16153
rect 8666 16079 8722 16088
rect 8680 15978 8708 16079
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8588 15830 8708 15858
rect 8482 15192 8538 15201
rect 8482 15127 8538 15136
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8206 13968 8262 13977
rect 8206 13903 8262 13912
rect 8312 13870 8340 14894
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8220 12782 8248 13738
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12986 8340 13126
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8312 12628 8340 12922
rect 8220 12600 8340 12628
rect 8114 11792 8170 11801
rect 8114 11727 8170 11736
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8128 11529 8156 11630
rect 8114 11520 8170 11529
rect 8114 11455 8170 11464
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7472 8502 7524 8508
rect 7654 8528 7710 8537
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7392 7478 7420 8434
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 6304 6868 7142
rect 6918 6760 6974 6769
rect 6918 6695 6974 6704
rect 7012 6724 7064 6730
rect 6932 6458 6960 6695
rect 7012 6666 7064 6672
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6920 6316 6972 6322
rect 6840 6276 6920 6304
rect 6840 5846 6868 6276
rect 6920 6258 6972 6264
rect 7024 6254 7052 6666
rect 7116 6322 7144 7346
rect 7286 6896 7342 6905
rect 7286 6831 7342 6840
rect 7194 6624 7250 6633
rect 7194 6559 7250 6568
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6748 3058 6776 3538
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6642 2952 6698 2961
rect 6840 2922 6868 4626
rect 6932 3194 6960 4966
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7024 2990 7052 3946
rect 7116 3602 7144 4082
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6642 2887 6698 2896
rect 6828 2916 6880 2922
rect 6828 2858 6880 2864
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6748 2378 6776 2790
rect 6840 2514 6868 2858
rect 6920 2848 6972 2854
rect 6918 2816 6920 2825
rect 6972 2816 6974 2825
rect 7116 2774 7144 3334
rect 6918 2751 6974 2760
rect 7024 2746 7144 2774
rect 7208 2774 7236 6559
rect 7300 5302 7328 6831
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7300 3602 7328 4150
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7286 3224 7342 3233
rect 7286 3159 7288 3168
rect 7340 3159 7342 3168
rect 7288 3130 7340 3136
rect 7208 2746 7328 2774
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 7024 2038 7052 2746
rect 7300 2666 7328 2746
rect 7116 2638 7328 2666
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 6552 1828 6604 1834
rect 6552 1770 6604 1776
rect 6276 1216 6328 1222
rect 6276 1158 6328 1164
rect 7116 800 7144 2638
rect 7392 1290 7420 7414
rect 7484 4593 7512 8502
rect 7654 8463 7710 8472
rect 7668 7993 7696 8463
rect 7654 7984 7710 7993
rect 7564 7948 7616 7954
rect 7654 7919 7710 7928
rect 7564 7890 7616 7896
rect 7576 7546 7604 7890
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7668 6798 7696 7482
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7576 5914 7604 6122
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7760 4706 7788 8774
rect 7576 4678 7788 4706
rect 7470 4584 7526 4593
rect 7470 4519 7526 4528
rect 7576 3058 7604 4678
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 3126 7696 3878
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7760 2009 7788 4490
rect 7852 3369 7880 8910
rect 7944 8498 7972 8910
rect 8036 8906 8064 9862
rect 8128 9602 8156 11222
rect 8220 10810 8248 12600
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8312 11665 8340 11698
rect 8298 11656 8354 11665
rect 8298 11591 8354 11600
rect 8298 11520 8354 11529
rect 8298 11455 8354 11464
rect 8312 11286 8340 11455
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8206 10704 8262 10713
rect 8206 10639 8262 10648
rect 8220 10062 8248 10639
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8312 9761 8340 11222
rect 8298 9752 8354 9761
rect 8298 9687 8354 9696
rect 8128 9574 8340 9602
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 8036 7721 8064 8842
rect 8128 8430 8156 9454
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8220 8974 8248 9114
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8022 7712 8078 7721
rect 8022 7647 8078 7656
rect 8036 6458 8064 7647
rect 8114 7576 8170 7585
rect 8114 7511 8170 7520
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8022 6352 8078 6361
rect 8022 6287 8078 6296
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4486 7972 4966
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7944 4146 7972 4422
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7930 4040 7986 4049
rect 7930 3975 7986 3984
rect 7838 3360 7894 3369
rect 7838 3295 7894 3304
rect 7852 2582 7880 3295
rect 7944 2990 7972 3975
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 8036 2774 8064 6287
rect 8128 5846 8156 7511
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8220 5030 8248 8910
rect 8312 6390 8340 9574
rect 8404 9178 8432 14962
rect 8496 14074 8524 15127
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8482 11928 8538 11937
rect 8482 11863 8538 11872
rect 8496 11626 8524 11863
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8482 11520 8538 11529
rect 8482 11455 8538 11464
rect 8496 11354 8524 11455
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8496 9450 8524 11086
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8588 8566 8616 14214
rect 8680 12730 8708 15830
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8772 13190 8800 14554
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8772 12850 8800 13126
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8680 12702 8800 12730
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8680 8378 8708 12038
rect 8772 9654 8800 12702
rect 8864 10810 8892 22510
rect 8956 22234 8984 23258
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 8956 14346 8984 22170
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8956 13938 8984 14282
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 12374 8984 12718
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8956 11150 8984 12174
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 9048 10674 9076 18566
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 9140 15745 9168 16118
rect 9232 16046 9260 25774
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9324 22778 9352 22918
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9324 16590 9352 22714
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9126 15736 9182 15745
rect 9126 15671 9182 15680
rect 9232 14550 9260 15982
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9140 11354 9168 12310
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8944 10532 8996 10538
rect 9128 10532 9180 10538
rect 8944 10474 8996 10480
rect 9048 10492 9128 10520
rect 8956 10266 8984 10474
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8588 8350 8708 8378
rect 8588 8106 8616 8350
rect 8588 8078 8708 8106
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8220 4214 8248 4694
rect 8312 4622 8340 5850
rect 8404 5778 8432 6666
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8496 4282 8524 7754
rect 8588 4865 8616 7822
rect 8574 4856 8630 4865
rect 8574 4791 8576 4800
rect 8628 4791 8630 4800
rect 8576 4762 8628 4768
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8128 3194 8156 4014
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8220 3058 8248 3674
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8036 2746 8340 2774
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 8312 2394 8340 2746
rect 8404 2514 8432 3470
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8588 2446 8616 4558
rect 8680 2774 8708 8078
rect 8772 3602 8800 9386
rect 8864 7954 8892 10066
rect 9048 9926 9076 10492
rect 9128 10474 9180 10480
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9126 9752 9182 9761
rect 9126 9687 9182 9696
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8956 9110 8984 9318
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 5914 8892 7890
rect 8956 7313 8984 8570
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8942 7304 8998 7313
rect 8942 7239 8998 7248
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8956 5234 8984 7239
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 9048 5030 9076 8026
rect 9140 7886 9168 9687
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7342 9168 7686
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9232 6497 9260 12582
rect 9416 12170 9444 26250
rect 11888 26240 11940 26246
rect 11888 26182 11940 26188
rect 10472 26140 10780 26149
rect 10472 26138 10478 26140
rect 10534 26138 10558 26140
rect 10614 26138 10638 26140
rect 10694 26138 10718 26140
rect 10774 26138 10780 26140
rect 10534 26086 10536 26138
rect 10716 26086 10718 26138
rect 10472 26084 10478 26086
rect 10534 26084 10558 26086
rect 10614 26084 10638 26086
rect 10694 26084 10718 26086
rect 10774 26084 10780 26086
rect 10472 26075 10780 26084
rect 10472 25052 10780 25061
rect 10472 25050 10478 25052
rect 10534 25050 10558 25052
rect 10614 25050 10638 25052
rect 10694 25050 10718 25052
rect 10774 25050 10780 25052
rect 10534 24998 10536 25050
rect 10716 24998 10718 25050
rect 10472 24996 10478 24998
rect 10534 24996 10558 24998
rect 10614 24996 10638 24998
rect 10694 24996 10718 24998
rect 10774 24996 10780 24998
rect 10472 24987 10780 24996
rect 10324 24132 10376 24138
rect 10324 24074 10376 24080
rect 10336 22710 10364 24074
rect 10472 23964 10780 23973
rect 10472 23962 10478 23964
rect 10534 23962 10558 23964
rect 10614 23962 10638 23964
rect 10694 23962 10718 23964
rect 10774 23962 10780 23964
rect 10534 23910 10536 23962
rect 10716 23910 10718 23962
rect 10472 23908 10478 23910
rect 10534 23908 10558 23910
rect 10614 23908 10638 23910
rect 10694 23908 10718 23910
rect 10774 23908 10780 23910
rect 10472 23899 10780 23908
rect 11060 23792 11112 23798
rect 11060 23734 11112 23740
rect 10472 22876 10780 22885
rect 10472 22874 10478 22876
rect 10534 22874 10558 22876
rect 10614 22874 10638 22876
rect 10694 22874 10718 22876
rect 10774 22874 10780 22876
rect 10534 22822 10536 22874
rect 10716 22822 10718 22874
rect 10472 22820 10478 22822
rect 10534 22820 10558 22822
rect 10614 22820 10638 22822
rect 10694 22820 10718 22822
rect 10774 22820 10780 22822
rect 10472 22811 10780 22820
rect 10324 22704 10376 22710
rect 10324 22646 10376 22652
rect 10472 21788 10780 21797
rect 10472 21786 10478 21788
rect 10534 21786 10558 21788
rect 10614 21786 10638 21788
rect 10694 21786 10718 21788
rect 10774 21786 10780 21788
rect 10534 21734 10536 21786
rect 10716 21734 10718 21786
rect 10472 21732 10478 21734
rect 10534 21732 10558 21734
rect 10614 21732 10638 21734
rect 10694 21732 10718 21734
rect 10774 21732 10780 21734
rect 10472 21723 10780 21732
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9508 14278 9536 17206
rect 9600 14482 9628 19450
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9692 15502 9720 16050
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9416 12073 9444 12106
rect 9402 12064 9458 12073
rect 9402 11999 9458 12008
rect 9508 11937 9536 14214
rect 9494 11928 9550 11937
rect 9312 11892 9364 11898
rect 9494 11863 9550 11872
rect 9312 11834 9364 11840
rect 9324 11014 9352 11834
rect 9600 11778 9628 14418
rect 9784 13394 9812 15506
rect 9876 14958 9904 20742
rect 10230 19408 10286 19417
rect 10230 19343 10286 19352
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9956 14544 10008 14550
rect 9956 14486 10008 14492
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9692 12850 9720 13262
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9692 12434 9720 12650
rect 9692 12406 9812 12434
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9508 11750 9628 11778
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 11218 9444 11494
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10810 9444 10826
rect 9324 10804 9456 10810
rect 9324 10798 9404 10804
rect 9324 10198 9352 10798
rect 9404 10746 9456 10752
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9324 9518 9352 9998
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9324 7342 9352 9454
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9218 6488 9274 6497
rect 9218 6423 9274 6432
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5545 9168 6258
rect 9324 6186 9352 6598
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9126 5536 9182 5545
rect 9126 5471 9182 5480
rect 9416 5370 9444 10610
rect 9508 8634 9536 11750
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 9738 9628 11562
rect 9692 10266 9720 12038
rect 9784 11898 9812 12406
rect 9876 12322 9904 13262
rect 9968 13258 9996 14486
rect 10060 14006 10088 15846
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 10152 12850 10180 15302
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9968 12442 9996 12786
rect 10244 12730 10272 19343
rect 10336 15162 10364 20810
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10472 20700 10780 20709
rect 10472 20698 10478 20700
rect 10534 20698 10558 20700
rect 10614 20698 10638 20700
rect 10694 20698 10718 20700
rect 10774 20698 10780 20700
rect 10534 20646 10536 20698
rect 10716 20646 10718 20698
rect 10472 20644 10478 20646
rect 10534 20644 10558 20646
rect 10614 20644 10638 20646
rect 10694 20644 10718 20646
rect 10774 20644 10780 20646
rect 10472 20635 10780 20644
rect 10472 19612 10780 19621
rect 10472 19610 10478 19612
rect 10534 19610 10558 19612
rect 10614 19610 10638 19612
rect 10694 19610 10718 19612
rect 10774 19610 10780 19612
rect 10534 19558 10536 19610
rect 10716 19558 10718 19610
rect 10472 19556 10478 19558
rect 10534 19556 10558 19558
rect 10614 19556 10638 19558
rect 10694 19556 10718 19558
rect 10774 19556 10780 19558
rect 10472 19547 10780 19556
rect 10472 18524 10780 18533
rect 10472 18522 10478 18524
rect 10534 18522 10558 18524
rect 10614 18522 10638 18524
rect 10694 18522 10718 18524
rect 10774 18522 10780 18524
rect 10534 18470 10536 18522
rect 10716 18470 10718 18522
rect 10472 18468 10478 18470
rect 10534 18468 10558 18470
rect 10614 18468 10638 18470
rect 10694 18468 10718 18470
rect 10774 18468 10780 18470
rect 10472 18459 10780 18468
rect 10472 17436 10780 17445
rect 10472 17434 10478 17436
rect 10534 17434 10558 17436
rect 10614 17434 10638 17436
rect 10694 17434 10718 17436
rect 10774 17434 10780 17436
rect 10534 17382 10536 17434
rect 10716 17382 10718 17434
rect 10472 17380 10478 17382
rect 10534 17380 10558 17382
rect 10614 17380 10638 17382
rect 10694 17380 10718 17382
rect 10774 17380 10780 17382
rect 10472 17371 10780 17380
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10472 16348 10780 16357
rect 10472 16346 10478 16348
rect 10534 16346 10558 16348
rect 10614 16346 10638 16348
rect 10694 16346 10718 16348
rect 10774 16346 10780 16348
rect 10534 16294 10536 16346
rect 10716 16294 10718 16346
rect 10472 16292 10478 16294
rect 10534 16292 10558 16294
rect 10614 16292 10638 16294
rect 10694 16292 10718 16294
rect 10774 16292 10780 16294
rect 10472 16283 10780 16292
rect 10472 15260 10780 15269
rect 10472 15258 10478 15260
rect 10534 15258 10558 15260
rect 10614 15258 10638 15260
rect 10694 15258 10718 15260
rect 10774 15258 10780 15260
rect 10534 15206 10536 15258
rect 10716 15206 10718 15258
rect 10472 15204 10478 15206
rect 10534 15204 10558 15206
rect 10614 15204 10638 15206
rect 10694 15204 10718 15206
rect 10774 15204 10780 15206
rect 10472 15195 10780 15204
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10336 14929 10364 15098
rect 10322 14920 10378 14929
rect 10322 14855 10378 14864
rect 10888 14657 10916 17070
rect 10980 16250 11008 20742
rect 11072 19281 11100 23734
rect 11520 23656 11572 23662
rect 11520 23598 11572 23604
rect 11244 23044 11296 23050
rect 11244 22986 11296 22992
rect 11256 22642 11284 22986
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11256 19854 11284 22578
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11348 20466 11376 22510
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11348 19378 11376 19994
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11058 19272 11114 19281
rect 11058 19207 11114 19216
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 11150 16552 11206 16561
rect 11150 16487 11206 16496
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11058 16008 11114 16017
rect 11058 15943 11060 15952
rect 11112 15943 11114 15952
rect 11060 15914 11112 15920
rect 11164 15094 11192 16487
rect 11256 15162 11284 18294
rect 11334 15328 11390 15337
rect 11334 15263 11390 15272
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 10874 14648 10930 14657
rect 10874 14583 10930 14592
rect 10876 14476 10928 14482
rect 10928 14436 11008 14464
rect 10876 14418 10928 14424
rect 10472 14172 10780 14181
rect 10472 14170 10478 14172
rect 10534 14170 10558 14172
rect 10614 14170 10638 14172
rect 10694 14170 10718 14172
rect 10774 14170 10780 14172
rect 10534 14118 10536 14170
rect 10716 14118 10718 14170
rect 10472 14116 10478 14118
rect 10534 14116 10558 14118
rect 10614 14116 10638 14118
rect 10694 14116 10718 14118
rect 10774 14116 10780 14118
rect 10472 14107 10780 14116
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10520 13802 10548 13874
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10060 12702 10272 12730
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9876 12294 9996 12322
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9876 11762 9904 12174
rect 9968 12170 9996 12294
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9954 12064 10010 12073
rect 9954 11999 10010 12008
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9876 11257 9904 11698
rect 9862 11248 9918 11257
rect 9862 11183 9918 11192
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9770 10160 9826 10169
rect 9770 10095 9826 10104
rect 9784 9976 9812 10095
rect 9864 9988 9916 9994
rect 9784 9948 9864 9976
rect 9864 9930 9916 9936
rect 9770 9888 9826 9897
rect 9770 9823 9826 9832
rect 9600 9710 9720 9738
rect 9692 9654 9720 9710
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9680 9512 9732 9518
rect 9784 9489 9812 9823
rect 9862 9752 9918 9761
rect 9862 9687 9918 9696
rect 9680 9454 9732 9460
rect 9770 9480 9826 9489
rect 9600 9178 9628 9454
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9692 9042 9720 9454
rect 9770 9415 9826 9424
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9770 8936 9826 8945
rect 9680 8900 9732 8906
rect 9770 8871 9826 8880
rect 9680 8842 9732 8848
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9692 8480 9720 8842
rect 9508 8452 9720 8480
rect 9508 6202 9536 8452
rect 9784 8430 9812 8871
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9876 8106 9904 9687
rect 9968 8294 9996 11999
rect 10060 10742 10088 12702
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9876 8078 9996 8106
rect 9862 7848 9918 7857
rect 9862 7783 9918 7792
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7206 9628 7686
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9586 6216 9642 6225
rect 9508 6174 9586 6202
rect 9586 6151 9642 6160
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9600 5234 9628 6151
rect 9678 5672 9734 5681
rect 9678 5607 9734 5616
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9232 4554 9260 4762
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8864 2990 8892 3878
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8680 2746 8984 2774
rect 8576 2440 8628 2446
rect 8312 2366 8432 2394
rect 8576 2382 8628 2388
rect 8956 2378 8984 2746
rect 9508 2582 9536 4966
rect 9692 4622 9720 5607
rect 9784 5574 9812 6734
rect 9876 6662 9904 7783
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9862 6488 9918 6497
rect 9862 6423 9918 6432
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9692 4486 9720 4558
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9692 3466 9720 4014
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 7746 2000 7802 2009
rect 7746 1935 7802 1944
rect 7380 1284 7432 1290
rect 7380 1226 7432 1232
rect 8404 800 8432 2366
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8496 1562 8524 2246
rect 9508 1902 9536 2518
rect 9784 2417 9812 4626
rect 9876 3126 9904 6423
rect 9968 5930 9996 8078
rect 10060 6361 10088 10202
rect 10152 8566 10180 12582
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10244 12345 10272 12378
rect 10230 12336 10286 12345
rect 10230 12271 10286 12280
rect 10232 12096 10284 12102
rect 10336 12073 10364 13738
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10472 13084 10780 13093
rect 10472 13082 10478 13084
rect 10534 13082 10558 13084
rect 10614 13082 10638 13084
rect 10694 13082 10718 13084
rect 10774 13082 10780 13084
rect 10534 13030 10536 13082
rect 10716 13030 10718 13082
rect 10472 13028 10478 13030
rect 10534 13028 10558 13030
rect 10614 13028 10638 13030
rect 10694 13028 10718 13030
rect 10774 13028 10780 13030
rect 10472 13019 10780 13028
rect 10888 12866 10916 13126
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10796 12838 10916 12866
rect 10520 12238 10548 12786
rect 10796 12646 10824 12838
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10612 12170 10640 12378
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10796 12102 10824 12310
rect 10784 12096 10836 12102
rect 10232 12038 10284 12044
rect 10322 12064 10378 12073
rect 10244 11121 10272 12038
rect 10784 12038 10836 12044
rect 10322 11999 10378 12008
rect 10472 11996 10780 12005
rect 10472 11994 10478 11996
rect 10534 11994 10558 11996
rect 10614 11994 10638 11996
rect 10694 11994 10718 11996
rect 10774 11994 10780 11996
rect 10534 11942 10536 11994
rect 10716 11942 10718 11994
rect 10472 11940 10478 11942
rect 10534 11940 10558 11942
rect 10614 11940 10638 11942
rect 10694 11940 10718 11942
rect 10774 11940 10780 11942
rect 10472 11931 10780 11940
rect 10784 11756 10836 11762
rect 10888 11744 10916 12718
rect 10980 11898 11008 14436
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 11072 12986 11100 13194
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11256 12374 11284 14758
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10836 11716 11008 11744
rect 10784 11698 10836 11704
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10230 11112 10286 11121
rect 10230 11047 10286 11056
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10674 10272 10950
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10244 10538 10272 10610
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10138 8392 10194 8401
rect 10138 8327 10194 8336
rect 10152 6798 10180 8327
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10046 6352 10102 6361
rect 10046 6287 10102 6296
rect 9968 5902 10088 5930
rect 10060 3602 10088 5902
rect 10152 5166 10180 6734
rect 10244 6458 10272 10202
rect 10336 9625 10364 11630
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10428 11336 10456 11562
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10508 11348 10560 11354
rect 10428 11308 10508 11336
rect 10508 11290 10560 11296
rect 10472 10908 10780 10917
rect 10472 10906 10478 10908
rect 10534 10906 10558 10908
rect 10614 10906 10638 10908
rect 10694 10906 10718 10908
rect 10774 10906 10780 10908
rect 10534 10854 10536 10906
rect 10716 10854 10718 10906
rect 10472 10852 10478 10854
rect 10534 10852 10558 10854
rect 10614 10852 10638 10854
rect 10694 10852 10718 10854
rect 10774 10852 10780 10854
rect 10472 10843 10780 10852
rect 10472 9820 10780 9829
rect 10472 9818 10478 9820
rect 10534 9818 10558 9820
rect 10614 9818 10638 9820
rect 10694 9818 10718 9820
rect 10774 9818 10780 9820
rect 10534 9766 10536 9818
rect 10716 9766 10718 9818
rect 10472 9764 10478 9766
rect 10534 9764 10558 9766
rect 10614 9764 10638 9766
rect 10694 9764 10718 9766
rect 10774 9764 10780 9766
rect 10472 9755 10780 9764
rect 10322 9616 10378 9625
rect 10322 9551 10378 9560
rect 10336 9042 10364 9551
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10414 9344 10470 9353
rect 10414 9279 10470 9288
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10428 8974 10456 9279
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10612 8906 10640 9386
rect 10782 9208 10838 9217
rect 10782 9143 10838 9152
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10796 8838 10824 9143
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10472 8732 10780 8741
rect 10472 8730 10478 8732
rect 10534 8730 10558 8732
rect 10614 8730 10638 8732
rect 10694 8730 10718 8732
rect 10774 8730 10780 8732
rect 10534 8678 10536 8730
rect 10716 8678 10718 8730
rect 10472 8676 10478 8678
rect 10534 8676 10558 8678
rect 10614 8676 10638 8678
rect 10694 8676 10718 8678
rect 10774 8676 10780 8678
rect 10472 8667 10780 8676
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10796 8401 10824 8502
rect 10782 8392 10838 8401
rect 10782 8327 10838 8336
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 8090 10824 8230
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10322 7984 10378 7993
rect 10322 7919 10378 7928
rect 10690 7984 10746 7993
rect 10690 7919 10692 7928
rect 10336 7177 10364 7919
rect 10744 7919 10746 7928
rect 10692 7890 10744 7896
rect 10472 7644 10780 7653
rect 10472 7642 10478 7644
rect 10534 7642 10558 7644
rect 10614 7642 10638 7644
rect 10694 7642 10718 7644
rect 10774 7642 10780 7644
rect 10534 7590 10536 7642
rect 10716 7590 10718 7642
rect 10472 7588 10478 7590
rect 10534 7588 10558 7590
rect 10614 7588 10638 7590
rect 10694 7588 10718 7590
rect 10774 7588 10780 7590
rect 10472 7579 10780 7588
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10322 7168 10378 7177
rect 10322 7103 10378 7112
rect 10428 6746 10456 7414
rect 10888 7410 10916 11494
rect 10980 9874 11008 11716
rect 11164 11257 11192 12038
rect 11256 11762 11284 12174
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11150 11248 11206 11257
rect 11150 11183 11206 11192
rect 11150 10704 11206 10713
rect 11060 10668 11112 10674
rect 11150 10639 11206 10648
rect 11060 10610 11112 10616
rect 11072 10198 11100 10610
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 11164 9994 11192 10639
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 10980 9846 11192 9874
rect 11058 9752 11114 9761
rect 11058 9687 11114 9696
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10980 7818 11008 8978
rect 11072 7954 11100 9687
rect 11164 9654 11192 9846
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11150 8664 11206 8673
rect 11150 8599 11206 8608
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10506 7168 10562 7177
rect 10506 7103 10562 7112
rect 10520 6866 10548 7103
rect 10874 6896 10930 6905
rect 10508 6860 10560 6866
rect 10980 6866 11008 7754
rect 10874 6831 10930 6840
rect 10968 6860 11020 6866
rect 10508 6802 10560 6808
rect 10336 6718 10456 6746
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10230 5808 10286 5817
rect 10230 5743 10286 5752
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10138 4176 10194 4185
rect 10244 4146 10272 5743
rect 10336 4321 10364 6718
rect 10472 6556 10780 6565
rect 10472 6554 10478 6556
rect 10534 6554 10558 6556
rect 10614 6554 10638 6556
rect 10694 6554 10718 6556
rect 10774 6554 10780 6556
rect 10534 6502 10536 6554
rect 10716 6502 10718 6554
rect 10472 6500 10478 6502
rect 10534 6500 10558 6502
rect 10614 6500 10638 6502
rect 10694 6500 10718 6502
rect 10774 6500 10780 6502
rect 10472 6491 10780 6500
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10506 6352 10562 6361
rect 10506 6287 10562 6296
rect 10520 6118 10548 6287
rect 10796 6118 10824 6394
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10888 5914 10916 6831
rect 10968 6802 11020 6808
rect 11058 6352 11114 6361
rect 10968 6316 11020 6322
rect 11058 6287 11114 6296
rect 10968 6258 11020 6264
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10472 5468 10780 5477
rect 10472 5466 10478 5468
rect 10534 5466 10558 5468
rect 10614 5466 10638 5468
rect 10694 5466 10718 5468
rect 10774 5466 10780 5468
rect 10534 5414 10536 5466
rect 10716 5414 10718 5466
rect 10472 5412 10478 5414
rect 10534 5412 10558 5414
rect 10614 5412 10638 5414
rect 10694 5412 10718 5414
rect 10774 5412 10780 5414
rect 10472 5403 10780 5412
rect 10980 5370 11008 6258
rect 11072 5778 11100 6287
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10874 4856 10930 4865
rect 10874 4791 10930 4800
rect 10888 4690 10916 4791
rect 10980 4690 11008 5306
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 11072 4826 11100 5238
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 11164 4622 11192 8599
rect 11256 8498 11284 11698
rect 11348 10062 11376 15263
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11440 12238 11468 15030
rect 11532 14958 11560 23598
rect 11900 23118 11928 26182
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 11992 23662 12020 24210
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11888 23112 11940 23118
rect 11888 23054 11940 23060
rect 11992 22094 12020 23598
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 11900 22066 12020 22094
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11624 14822 11652 19790
rect 11716 16250 11744 21898
rect 11900 17134 11928 22066
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11992 20602 12020 21626
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11808 16114 11836 16594
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11716 15162 11744 15642
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11808 15026 11836 16050
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11900 15706 11928 15846
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11900 15162 11928 15302
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11992 15094 12020 20334
rect 12070 15192 12126 15201
rect 12070 15127 12126 15136
rect 11980 15088 12032 15094
rect 11886 15056 11942 15065
rect 11796 15020 11848 15026
rect 11980 15030 12032 15036
rect 12084 15026 12112 15127
rect 12176 15065 12204 23462
rect 12268 19378 12296 24754
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12268 18766 12296 19314
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12268 16658 12296 18702
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 12268 15162 12296 16458
rect 12360 15434 12388 23802
rect 12452 23322 12480 24346
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12452 19378 12480 22034
rect 12544 21146 12572 22578
rect 12636 21554 12664 24006
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12636 21350 12664 21490
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12532 21140 12584 21146
rect 12532 21082 12584 21088
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12532 20936 12584 20942
rect 12636 20913 12664 20946
rect 12532 20878 12584 20884
rect 12622 20904 12678 20913
rect 12544 20534 12572 20878
rect 12622 20839 12678 20848
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 12544 19854 12572 20470
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18290 12480 19314
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12438 15736 12494 15745
rect 12438 15671 12494 15680
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12162 15056 12218 15065
rect 11886 14991 11942 15000
rect 12072 15020 12124 15026
rect 11796 14962 11848 14968
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11794 14648 11850 14657
rect 11794 14583 11850 14592
rect 11808 14414 11836 14583
rect 11900 14414 11928 14991
rect 12162 14991 12218 15000
rect 12072 14962 12124 14968
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 12084 14346 12112 14962
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11624 13433 11652 14010
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11610 13424 11666 13433
rect 11610 13359 11666 13368
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11242 8120 11298 8129
rect 11242 8055 11298 8064
rect 11256 7585 11284 8055
rect 11242 7576 11298 7585
rect 11242 7511 11298 7520
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11256 6730 11284 7278
rect 11348 6730 11376 8978
rect 11440 8634 11468 10406
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11256 4622 11284 6258
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11348 5166 11376 5646
rect 11440 5574 11468 8434
rect 11532 7818 11560 12650
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11624 11354 11652 12038
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11716 10826 11744 12038
rect 11794 11384 11850 11393
rect 11794 11319 11850 11328
rect 11808 11150 11836 11319
rect 11900 11218 11928 12174
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11992 11150 12020 13874
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 13258 12112 13670
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12084 12753 12112 12786
rect 12070 12744 12126 12753
rect 12070 12679 12126 12688
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11624 10798 11744 10826
rect 11624 9518 11652 10798
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11716 9382 11744 10610
rect 11794 10296 11850 10305
rect 11794 10231 11850 10240
rect 11808 9761 11836 10231
rect 11900 9994 11928 10950
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11794 9752 11850 9761
rect 11794 9687 11850 9696
rect 11886 9616 11942 9625
rect 11992 9586 12020 11086
rect 12070 10976 12126 10985
rect 12070 10911 12126 10920
rect 12084 10742 12112 10911
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 12084 9897 12112 10406
rect 12070 9888 12126 9897
rect 12070 9823 12126 9832
rect 11886 9551 11942 9560
rect 11980 9580 12032 9586
rect 11900 9518 11928 9551
rect 11980 9522 12032 9528
rect 11888 9512 11940 9518
rect 11794 9480 11850 9489
rect 11888 9454 11940 9460
rect 11794 9415 11850 9424
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11808 8888 11836 9415
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9081 11928 9318
rect 11886 9072 11942 9081
rect 11886 9007 11942 9016
rect 11888 8900 11940 8906
rect 11808 8860 11888 8888
rect 11888 8842 11940 8848
rect 11992 8786 12020 9522
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 11808 8758 12020 8786
rect 11610 8256 11666 8265
rect 11610 8191 11666 8200
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11624 5953 11652 8191
rect 11808 7410 11836 8758
rect 12084 8566 12112 9386
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11716 7002 11744 7142
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11610 5944 11666 5953
rect 11610 5879 11666 5888
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11256 4468 11284 4558
rect 11164 4440 11284 4468
rect 10472 4380 10780 4389
rect 10472 4378 10478 4380
rect 10534 4378 10558 4380
rect 10614 4378 10638 4380
rect 10694 4378 10718 4380
rect 10774 4378 10780 4380
rect 10534 4326 10536 4378
rect 10716 4326 10718 4378
rect 10472 4324 10478 4326
rect 10534 4324 10558 4326
rect 10614 4324 10638 4326
rect 10694 4324 10718 4326
rect 10774 4324 10780 4326
rect 10322 4312 10378 4321
rect 10472 4315 10780 4324
rect 10322 4247 10378 4256
rect 10336 4214 10364 4247
rect 10324 4208 10376 4214
rect 10692 4208 10744 4214
rect 10324 4150 10376 4156
rect 10690 4176 10692 4185
rect 10744 4176 10746 4185
rect 10138 4111 10194 4120
rect 10232 4140 10284 4146
rect 10152 4078 10180 4111
rect 10690 4111 10746 4120
rect 10232 4082 10284 4088
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3602 10180 3878
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 10060 2446 10088 3538
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10472 3292 10780 3301
rect 10472 3290 10478 3292
rect 10534 3290 10558 3292
rect 10614 3290 10638 3292
rect 10694 3290 10718 3292
rect 10774 3290 10780 3292
rect 10534 3238 10536 3290
rect 10716 3238 10718 3290
rect 10472 3236 10478 3238
rect 10534 3236 10558 3238
rect 10614 3236 10638 3238
rect 10694 3236 10718 3238
rect 10774 3236 10780 3238
rect 10472 3227 10780 3236
rect 11072 3233 11100 3470
rect 11058 3224 11114 3233
rect 11058 3159 11114 3168
rect 11164 3108 11192 4440
rect 11242 3632 11298 3641
rect 11242 3567 11298 3576
rect 11256 3126 11284 3567
rect 11348 3534 11376 5102
rect 11808 3942 11836 5578
rect 11900 5302 11928 8434
rect 12176 8378 12204 12786
rect 12268 12714 12296 14282
rect 12360 14113 12388 14894
rect 12452 14385 12480 15671
rect 12438 14376 12494 14385
rect 12438 14311 12494 14320
rect 12346 14104 12402 14113
rect 12346 14039 12402 14048
rect 12544 13802 12572 16730
rect 12636 16182 12664 20470
rect 12728 19310 12756 24550
rect 13004 23730 13032 25842
rect 13096 24750 13124 26386
rect 14936 26382 14964 28478
rect 16118 28354 16174 29154
rect 18050 28506 18106 29154
rect 19982 28506 20038 29154
rect 21914 28506 21970 29154
rect 23202 28506 23258 29154
rect 18050 28478 18184 28506
rect 18050 28354 18106 28478
rect 16132 28286 16160 28354
rect 16120 28280 16172 28286
rect 16120 28222 16172 28228
rect 17132 28280 17184 28286
rect 17132 28222 17184 28228
rect 15233 26684 15541 26693
rect 15233 26682 15239 26684
rect 15295 26682 15319 26684
rect 15375 26682 15399 26684
rect 15455 26682 15479 26684
rect 15535 26682 15541 26684
rect 15295 26630 15297 26682
rect 15477 26630 15479 26682
rect 15233 26628 15239 26630
rect 15295 26628 15319 26630
rect 15375 26628 15399 26630
rect 15455 26628 15479 26630
rect 15535 26628 15541 26630
rect 15233 26619 15541 26628
rect 15568 26512 15620 26518
rect 15568 26454 15620 26460
rect 16120 26512 16172 26518
rect 16120 26454 16172 26460
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 14924 26240 14976 26246
rect 14924 26182 14976 26188
rect 14832 25764 14884 25770
rect 14832 25706 14884 25712
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13556 24750 13584 25094
rect 13084 24744 13136 24750
rect 13082 24712 13084 24721
rect 13544 24744 13596 24750
rect 13136 24712 13138 24721
rect 13544 24686 13596 24692
rect 13082 24647 13138 24656
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13464 22982 13492 24006
rect 13556 23594 13584 24686
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13544 23588 13596 23594
rect 13544 23530 13596 23536
rect 13556 23186 13584 23530
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13740 23118 13768 23666
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13544 23044 13596 23050
rect 13544 22986 13596 22992
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 12808 21888 12860 21894
rect 12992 21888 13044 21894
rect 12860 21836 12992 21842
rect 12808 21830 13044 21836
rect 12820 21814 13032 21830
rect 13096 21570 13124 22510
rect 12820 21554 13124 21570
rect 12808 21548 13124 21554
rect 12860 21542 13124 21548
rect 12808 21490 12860 21496
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 12820 20330 12848 21082
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12992 20868 13044 20874
rect 12992 20810 13044 20816
rect 12912 20534 12940 20810
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 13004 20262 13032 20810
rect 13096 20262 13124 21542
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 12900 19848 12952 19854
rect 13004 19836 13032 20198
rect 12952 19808 13032 19836
rect 12900 19790 12952 19796
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12728 16250 12756 16390
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12728 15745 12756 15914
rect 12714 15736 12770 15745
rect 12714 15671 12770 15680
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12636 15366 12664 15506
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 13938 12664 15302
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12728 14482 12756 14894
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12360 13190 12388 13330
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12753 12480 13126
rect 12438 12744 12494 12753
rect 12256 12708 12308 12714
rect 12438 12679 12494 12688
rect 12256 12650 12308 12656
rect 12544 12646 12572 13738
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 11992 8350 12204 8378
rect 11992 5846 12020 8350
rect 12070 7984 12126 7993
rect 12070 7919 12126 7928
rect 12084 7274 12112 7919
rect 12268 7721 12296 11494
rect 12360 8106 12388 12582
rect 12544 12442 12572 12582
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12636 11762 12664 13874
rect 12714 12744 12770 12753
rect 12714 12679 12770 12688
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 12452 11354 12480 11562
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12452 8514 12480 11290
rect 12636 11218 12664 11698
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12624 10600 12676 10606
rect 12728 10554 12756 12679
rect 12676 10548 12756 10554
rect 12624 10542 12756 10548
rect 12636 10526 12756 10542
rect 12530 10024 12586 10033
rect 12530 9959 12586 9968
rect 12544 9926 12572 9959
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12728 9654 12756 10526
rect 12820 10130 12848 19654
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12912 15978 12940 16458
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12912 12850 12940 15506
rect 13004 14346 13032 19382
rect 13096 14906 13124 20198
rect 13188 20058 13216 21490
rect 13280 21486 13308 22918
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13280 20398 13308 20878
rect 13268 20392 13320 20398
rect 13268 20334 13320 20340
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13280 19854 13308 20334
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13188 17202 13216 18226
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13188 16114 13216 17138
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13266 15056 13322 15065
rect 13266 14991 13322 15000
rect 13096 14878 13216 14906
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14414 13124 14758
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13004 13138 13032 14282
rect 13188 13410 13216 14878
rect 13280 14550 13308 14991
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13268 14408 13320 14414
rect 13266 14376 13268 14385
rect 13320 14376 13322 14385
rect 13266 14311 13322 14320
rect 13188 13394 13308 13410
rect 13372 13394 13400 21830
rect 13464 20806 13492 22918
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13450 19544 13506 19553
rect 13450 19479 13506 19488
rect 13464 14550 13492 19479
rect 13556 16182 13584 22986
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13648 21010 13676 22102
rect 13728 21956 13780 21962
rect 13728 21898 13780 21904
rect 13740 21078 13768 21898
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13726 20360 13782 20369
rect 13726 20295 13728 20304
rect 13780 20295 13782 20304
rect 13728 20266 13780 20272
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13648 19689 13676 19722
rect 13634 19680 13690 19689
rect 13634 19615 13690 19624
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13648 16590 13676 17274
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13740 15706 13768 19450
rect 13832 19378 13860 25638
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13924 22642 13952 25230
rect 14844 25226 14872 25706
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14096 24880 14148 24886
rect 14096 24822 14148 24828
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13924 22030 13952 22578
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13832 16658 13860 16730
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13818 16280 13874 16289
rect 13818 16215 13874 16224
rect 13832 16017 13860 16215
rect 13818 16008 13874 16017
rect 13818 15943 13874 15952
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13648 15416 13676 15642
rect 13648 15388 13768 15416
rect 13740 15026 13768 15388
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13464 14249 13492 14282
rect 13450 14240 13506 14249
rect 13450 14175 13506 14184
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13188 13388 13320 13394
rect 13188 13382 13268 13388
rect 13268 13330 13320 13336
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13176 13320 13228 13326
rect 13174 13288 13176 13297
rect 13228 13288 13230 13297
rect 13280 13258 13308 13330
rect 13174 13223 13230 13232
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13004 13110 13400 13138
rect 13176 12912 13228 12918
rect 13268 12912 13320 12918
rect 13176 12854 13228 12860
rect 13266 12880 13268 12889
rect 13320 12880 13322 12889
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 13188 12753 13216 12854
rect 13266 12815 13322 12824
rect 13174 12744 13230 12753
rect 13174 12679 13230 12688
rect 13280 12170 13308 12815
rect 13372 12238 13400 13110
rect 13464 12481 13492 13806
rect 13556 12986 13584 14826
rect 13818 14512 13874 14521
rect 13818 14447 13874 14456
rect 13832 13852 13860 14447
rect 13924 14414 13952 19994
rect 14016 19514 14044 23666
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14108 19417 14136 24822
rect 14844 24818 14872 25162
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14094 19408 14150 19417
rect 14094 19343 14150 19352
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 17202 14136 17614
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13832 13824 13952 13852
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13450 12472 13506 12481
rect 13450 12407 13506 12416
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13464 12084 13492 12407
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13372 12056 13492 12084
rect 13176 11824 13228 11830
rect 13174 11792 13176 11801
rect 13228 11792 13230 11801
rect 13174 11727 13230 11736
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12898 10296 12954 10305
rect 12898 10231 12954 10240
rect 12912 10198 12940 10231
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12716 9648 12768 9654
rect 12530 9616 12586 9625
rect 12716 9590 12768 9596
rect 12530 9551 12532 9560
rect 12584 9551 12586 9560
rect 12532 9522 12584 9528
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12530 9208 12586 9217
rect 12530 9143 12586 9152
rect 12544 9110 12572 9143
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12544 8634 12572 9046
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12452 8486 12572 8514
rect 12360 8078 12480 8106
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 12254 7712 12310 7721
rect 12254 7647 12310 7656
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12084 6186 12112 6938
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11992 5658 12020 5782
rect 11992 5630 12204 5658
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11992 4826 12020 5102
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 12084 4146 12112 5510
rect 12176 4486 12204 5630
rect 12268 4865 12296 7210
rect 12254 4856 12310 4865
rect 12254 4791 12310 4800
rect 12268 4690 12296 4791
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12360 4146 12388 7958
rect 12452 7188 12480 8078
rect 12544 7342 12572 8486
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12636 7256 12664 8434
rect 12728 7478 12756 9386
rect 12820 7954 12848 10066
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 8906 12940 9862
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12636 7228 12756 7256
rect 12452 7160 12664 7188
rect 12438 7032 12494 7041
rect 12438 6967 12494 6976
rect 12452 6798 12480 6967
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12530 6760 12586 6769
rect 12530 6695 12586 6704
rect 12544 6458 12572 6695
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12544 6225 12572 6394
rect 12530 6216 12586 6225
rect 12530 6151 12586 6160
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12254 4040 12310 4049
rect 12254 3975 12310 3984
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11348 3126 11376 3470
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11624 3194 11652 3402
rect 12176 3194 12204 3674
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 11072 3080 11192 3108
rect 11244 3120 11296 3126
rect 11072 2854 11100 3080
rect 11244 3062 11296 3068
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10048 2440 10100 2446
rect 9770 2408 9826 2417
rect 10048 2382 10100 2388
rect 9770 2343 9826 2352
rect 10472 2204 10780 2213
rect 10472 2202 10478 2204
rect 10534 2202 10558 2204
rect 10614 2202 10638 2204
rect 10694 2202 10718 2204
rect 10774 2202 10780 2204
rect 10534 2150 10536 2202
rect 10716 2150 10718 2202
rect 10472 2148 10478 2150
rect 10534 2148 10558 2150
rect 10614 2148 10638 2150
rect 10694 2148 10718 2150
rect 10774 2148 10780 2150
rect 10472 2139 10780 2148
rect 9496 1896 9548 1902
rect 9496 1838 9548 1844
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 11164 950 11192 2858
rect 12176 2774 12204 3130
rect 12084 2746 12204 2774
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11888 2576 11940 2582
rect 11888 2518 11940 2524
rect 11808 1154 11836 2518
rect 11900 2446 11928 2518
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 12084 2378 12112 2746
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12176 1970 12204 2246
rect 12164 1964 12216 1970
rect 12164 1906 12216 1912
rect 12176 1766 12204 1906
rect 12164 1760 12216 1766
rect 12164 1702 12216 1708
rect 11796 1148 11848 1154
rect 11796 1090 11848 1096
rect 11152 944 11204 950
rect 10244 870 10364 898
rect 11152 886 11204 892
rect 5540 128 5592 134
rect 5540 70 5592 76
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 10244 134 10272 870
rect 10336 800 10364 870
rect 12268 800 12296 3975
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 2038 12388 3538
rect 12452 2990 12480 4626
rect 12636 3466 12664 7160
rect 12728 6322 12756 7228
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12820 4010 12848 7346
rect 12912 6934 12940 8842
rect 13004 7478 13032 11494
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13004 5914 13032 6734
rect 13096 6254 13124 10134
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 9217 13216 9454
rect 13174 9208 13230 9217
rect 13174 9143 13230 9152
rect 13174 8800 13230 8809
rect 13174 8735 13230 8744
rect 13188 8566 13216 8735
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13188 7750 13216 8366
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13188 6089 13216 7346
rect 13174 6080 13230 6089
rect 13174 6015 13230 6024
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13280 5817 13308 8230
rect 13372 6390 13400 12056
rect 13556 11937 13584 12174
rect 13648 12170 13676 13262
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13740 12442 13768 12718
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13542 11928 13598 11937
rect 13542 11863 13598 11872
rect 13740 11558 13768 12106
rect 13832 11898 13860 12786
rect 13924 12102 13952 13824
rect 14016 12238 14044 15846
rect 14108 15570 14136 17138
rect 14200 16182 14228 24550
rect 14752 24274 14780 24686
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 14648 24064 14700 24070
rect 14648 24006 14700 24012
rect 14292 22710 14320 24006
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14292 19514 14320 19654
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14278 19408 14334 19417
rect 14278 19343 14334 19352
rect 14292 19242 14320 19343
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14188 16176 14240 16182
rect 14188 16118 14240 16124
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14108 15094 14136 15506
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 13977 14136 14350
rect 14094 13968 14150 13977
rect 14094 13903 14150 13912
rect 14200 12288 14228 15642
rect 14384 15502 14412 22918
rect 14660 22574 14688 24006
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14556 22432 14608 22438
rect 14752 22386 14780 24210
rect 14936 24206 14964 26182
rect 15233 25596 15541 25605
rect 15233 25594 15239 25596
rect 15295 25594 15319 25596
rect 15375 25594 15399 25596
rect 15455 25594 15479 25596
rect 15535 25594 15541 25596
rect 15295 25542 15297 25594
rect 15477 25542 15479 25594
rect 15233 25540 15239 25542
rect 15295 25540 15319 25542
rect 15375 25540 15399 25542
rect 15455 25540 15479 25542
rect 15535 25540 15541 25542
rect 15233 25531 15541 25540
rect 15233 24508 15541 24517
rect 15233 24506 15239 24508
rect 15295 24506 15319 24508
rect 15375 24506 15399 24508
rect 15455 24506 15479 24508
rect 15535 24506 15541 24508
rect 15295 24454 15297 24506
rect 15477 24454 15479 24506
rect 15233 24452 15239 24454
rect 15295 24452 15319 24454
rect 15375 24452 15399 24454
rect 15455 24452 15479 24454
rect 15535 24452 15541 24454
rect 15233 24443 15541 24452
rect 15016 24336 15068 24342
rect 15016 24278 15068 24284
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14556 22374 14608 22380
rect 14568 22094 14596 22374
rect 14476 22066 14596 22094
rect 14660 22358 14780 22386
rect 14476 20058 14504 22066
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14556 19984 14608 19990
rect 14556 19926 14608 19932
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14292 15144 14320 15370
rect 14292 15116 14412 15144
rect 14278 15056 14334 15065
rect 14278 14991 14334 15000
rect 14292 13530 14320 14991
rect 14384 14958 14412 15116
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14384 14260 14412 14894
rect 14476 14414 14504 19858
rect 14568 16522 14596 19926
rect 14556 16516 14608 16522
rect 14556 16458 14608 16464
rect 14554 15736 14610 15745
rect 14554 15671 14610 15680
rect 14568 14618 14596 15671
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14384 14232 14504 14260
rect 14476 14006 14504 14232
rect 14568 14074 14596 14554
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14108 12260 14228 12288
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13450 10840 13506 10849
rect 13450 10775 13506 10784
rect 13464 10742 13492 10775
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 9994 13492 10542
rect 13556 9994 13584 11086
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13450 9208 13506 9217
rect 13450 9143 13506 9152
rect 13464 9042 13492 9143
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13464 7342 13492 8978
rect 13648 8838 13676 11222
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 7886 13676 8774
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13648 6934 13676 7822
rect 13740 7410 13768 10406
rect 13924 9926 13952 11834
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 13740 6882 13768 7346
rect 13832 7206 13860 9658
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13924 9353 13952 9522
rect 13910 9344 13966 9353
rect 13910 9279 13966 9288
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13924 8634 13952 8978
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13740 6866 13860 6882
rect 13728 6860 13860 6866
rect 13780 6854 13860 6860
rect 13728 6802 13780 6808
rect 13542 6488 13598 6497
rect 13542 6423 13544 6432
rect 13596 6423 13598 6432
rect 13544 6394 13596 6400
rect 13832 6390 13860 6854
rect 14016 6798 14044 12174
rect 14108 10266 14136 12260
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13266 5808 13322 5817
rect 13266 5743 13322 5752
rect 13372 5302 13400 6054
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12912 2650 12940 4082
rect 13004 4078 13032 4558
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4185 13216 4422
rect 13174 4176 13230 4185
rect 13084 4140 13136 4146
rect 13174 4111 13230 4120
rect 13084 4082 13136 4088
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 3058 13032 3470
rect 13096 3398 13124 4082
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13096 3194 13124 3334
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13004 2582 13032 2994
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 13004 2360 13032 2518
rect 13176 2372 13228 2378
rect 13004 2332 13176 2360
rect 13176 2314 13228 2320
rect 12348 2032 12400 2038
rect 12348 1974 12400 1980
rect 13280 1737 13308 5238
rect 13358 4856 13414 4865
rect 13358 4791 13414 4800
rect 13372 4690 13400 4791
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 13372 3194 13400 4218
rect 13464 4214 13492 4626
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 13450 3496 13506 3505
rect 13450 3431 13506 3440
rect 13464 3233 13492 3431
rect 13450 3224 13506 3233
rect 13360 3188 13412 3194
rect 13450 3159 13506 3168
rect 13360 3130 13412 3136
rect 13556 1902 13584 5578
rect 13648 5574 13676 6054
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13648 2145 13676 3878
rect 13740 2774 13768 5850
rect 13924 5030 13952 6190
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 14016 4706 14044 6734
rect 14108 5710 14136 10202
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14096 5704 14148 5710
rect 14200 5692 14228 8978
rect 14292 8974 14320 13194
rect 14384 10266 14412 13942
rect 14568 13682 14596 14010
rect 14660 13938 14688 22358
rect 14844 22030 14872 23054
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 14936 20602 14964 24142
rect 15028 23798 15056 24278
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15212 24070 15240 24142
rect 15108 24064 15160 24070
rect 15108 24006 15160 24012
rect 15200 24064 15252 24070
rect 15200 24006 15252 24012
rect 15016 23792 15068 23798
rect 15016 23734 15068 23740
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14844 19378 14872 19994
rect 14936 19718 14964 20198
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 14936 19446 14964 19654
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14660 13734 14688 13874
rect 14476 13654 14596 13682
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14476 12889 14504 13654
rect 14646 13560 14702 13569
rect 14556 13524 14608 13530
rect 14752 13530 14780 18158
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 14414 14872 15302
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14646 13495 14702 13504
rect 14740 13524 14792 13530
rect 14556 13466 14608 13472
rect 14462 12880 14518 12889
rect 14462 12815 14518 12824
rect 14462 12336 14518 12345
rect 14462 12271 14518 12280
rect 14476 11558 14504 12271
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14462 10840 14518 10849
rect 14462 10775 14464 10784
rect 14516 10775 14518 10784
rect 14464 10746 14516 10752
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14476 9674 14504 10542
rect 14384 9646 14504 9674
rect 14384 9489 14412 9646
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14370 9480 14426 9489
rect 14370 9415 14426 9424
rect 14476 9110 14504 9522
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14384 8514 14412 8910
rect 14292 8362 14320 8502
rect 14384 8486 14432 8514
rect 14280 8356 14332 8362
rect 14404 8344 14432 8486
rect 14568 8430 14596 13466
rect 14660 12986 14688 13495
rect 14740 13466 14792 13472
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14660 9586 14688 12650
rect 14752 12238 14780 13126
rect 14844 12238 14872 13806
rect 14936 13326 14964 18022
rect 15028 16046 15056 21422
rect 15120 18193 15148 24006
rect 15580 23866 15608 26454
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 15568 23860 15620 23866
rect 15620 23820 15700 23848
rect 15568 23802 15620 23808
rect 15233 23420 15541 23429
rect 15233 23418 15239 23420
rect 15295 23418 15319 23420
rect 15375 23418 15399 23420
rect 15455 23418 15479 23420
rect 15535 23418 15541 23420
rect 15295 23366 15297 23418
rect 15477 23366 15479 23418
rect 15233 23364 15239 23366
rect 15295 23364 15319 23366
rect 15375 23364 15399 23366
rect 15455 23364 15479 23366
rect 15535 23364 15541 23366
rect 15233 23355 15541 23364
rect 15568 22704 15620 22710
rect 15568 22646 15620 22652
rect 15233 22332 15541 22341
rect 15233 22330 15239 22332
rect 15295 22330 15319 22332
rect 15375 22330 15399 22332
rect 15455 22330 15479 22332
rect 15535 22330 15541 22332
rect 15295 22278 15297 22330
rect 15477 22278 15479 22330
rect 15233 22276 15239 22278
rect 15295 22276 15319 22278
rect 15375 22276 15399 22278
rect 15455 22276 15479 22278
rect 15535 22276 15541 22278
rect 15233 22267 15541 22276
rect 15580 22098 15608 22646
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15233 21244 15541 21253
rect 15233 21242 15239 21244
rect 15295 21242 15319 21244
rect 15375 21242 15399 21244
rect 15455 21242 15479 21244
rect 15535 21242 15541 21244
rect 15295 21190 15297 21242
rect 15477 21190 15479 21242
rect 15233 21188 15239 21190
rect 15295 21188 15319 21190
rect 15375 21188 15399 21190
rect 15455 21188 15479 21190
rect 15535 21188 15541 21190
rect 15233 21179 15541 21188
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15233 20156 15541 20165
rect 15233 20154 15239 20156
rect 15295 20154 15319 20156
rect 15375 20154 15399 20156
rect 15455 20154 15479 20156
rect 15535 20154 15541 20156
rect 15295 20102 15297 20154
rect 15477 20102 15479 20154
rect 15233 20100 15239 20102
rect 15295 20100 15319 20102
rect 15375 20100 15399 20102
rect 15455 20100 15479 20102
rect 15535 20100 15541 20102
rect 15233 20091 15541 20100
rect 15233 19068 15541 19077
rect 15233 19066 15239 19068
rect 15295 19066 15319 19068
rect 15375 19066 15399 19068
rect 15455 19066 15479 19068
rect 15535 19066 15541 19068
rect 15295 19014 15297 19066
rect 15477 19014 15479 19066
rect 15233 19012 15239 19014
rect 15295 19012 15319 19014
rect 15375 19012 15399 19014
rect 15455 19012 15479 19014
rect 15535 19012 15541 19014
rect 15233 19003 15541 19012
rect 15106 18184 15162 18193
rect 15106 18119 15162 18128
rect 15233 17980 15541 17989
rect 15233 17978 15239 17980
rect 15295 17978 15319 17980
rect 15375 17978 15399 17980
rect 15455 17978 15479 17980
rect 15535 17978 15541 17980
rect 15295 17926 15297 17978
rect 15477 17926 15479 17978
rect 15233 17924 15239 17926
rect 15295 17924 15319 17926
rect 15375 17924 15399 17926
rect 15455 17924 15479 17926
rect 15535 17924 15541 17926
rect 15233 17915 15541 17924
rect 15233 16892 15541 16901
rect 15233 16890 15239 16892
rect 15295 16890 15319 16892
rect 15375 16890 15399 16892
rect 15455 16890 15479 16892
rect 15535 16890 15541 16892
rect 15295 16838 15297 16890
rect 15477 16838 15479 16890
rect 15233 16836 15239 16838
rect 15295 16836 15319 16838
rect 15375 16836 15399 16838
rect 15455 16836 15479 16838
rect 15535 16836 15541 16838
rect 15233 16827 15541 16836
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15120 16182 15148 16526
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15120 15706 15148 16118
rect 15396 16114 15424 16662
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 15198 16008 15254 16017
rect 15198 15943 15200 15952
rect 15252 15943 15254 15952
rect 15200 15914 15252 15920
rect 15233 15804 15541 15813
rect 15233 15802 15239 15804
rect 15295 15802 15319 15804
rect 15375 15802 15399 15804
rect 15455 15802 15479 15804
rect 15535 15802 15541 15804
rect 15295 15750 15297 15802
rect 15477 15750 15479 15802
rect 15233 15748 15239 15750
rect 15295 15748 15319 15750
rect 15375 15748 15399 15750
rect 15455 15748 15479 15750
rect 15535 15748 15541 15750
rect 15233 15739 15541 15748
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15028 14414 15056 15370
rect 15580 15201 15608 20538
rect 15672 18737 15700 23820
rect 15856 21690 15884 24142
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 16040 19553 16068 24142
rect 16026 19544 16082 19553
rect 16026 19479 16082 19488
rect 15658 18728 15714 18737
rect 15658 18663 15714 18672
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15672 17202 15700 17614
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15566 15192 15622 15201
rect 15566 15127 15622 15136
rect 15233 14716 15541 14725
rect 15233 14714 15239 14716
rect 15295 14714 15319 14716
rect 15375 14714 15399 14716
rect 15455 14714 15479 14716
rect 15535 14714 15541 14716
rect 15295 14662 15297 14714
rect 15477 14662 15479 14714
rect 15233 14660 15239 14662
rect 15295 14660 15319 14662
rect 15375 14660 15399 14662
rect 15455 14660 15479 14662
rect 15535 14660 15541 14662
rect 15106 14648 15162 14657
rect 15233 14651 15541 14660
rect 15106 14583 15162 14592
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14936 13190 14964 13262
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14740 12096 14792 12102
rect 14936 12084 14964 12922
rect 14740 12038 14792 12044
rect 14844 12056 14964 12084
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14280 8298 14332 8304
rect 14384 8316 14432 8344
rect 14384 8242 14412 8316
rect 14660 8294 14688 9522
rect 14752 9178 14780 12038
rect 14844 10062 14872 12056
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14936 10130 14964 10746
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 15028 9674 15056 14010
rect 15120 14006 15148 14583
rect 15672 14346 15700 16458
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15580 13870 15608 13942
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15120 13376 15148 13670
rect 15233 13628 15541 13637
rect 15233 13626 15239 13628
rect 15295 13626 15319 13628
rect 15375 13626 15399 13628
rect 15455 13626 15479 13628
rect 15535 13626 15541 13628
rect 15295 13574 15297 13626
rect 15477 13574 15479 13626
rect 15233 13572 15239 13574
rect 15295 13572 15319 13574
rect 15375 13572 15399 13574
rect 15455 13572 15479 13574
rect 15535 13572 15541 13574
rect 15233 13563 15541 13572
rect 15200 13388 15252 13394
rect 15120 13348 15200 13376
rect 15200 13330 15252 13336
rect 15580 13274 15608 13806
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15212 13246 15608 13274
rect 15672 13258 15700 13670
rect 15764 13326 15792 15982
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15660 13252 15712 13258
rect 15212 12986 15240 13246
rect 15660 13194 15712 13200
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15120 12753 15148 12786
rect 15106 12744 15162 12753
rect 15106 12679 15162 12688
rect 15304 12628 15332 13126
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 14844 9646 15056 9674
rect 15120 12600 15332 12628
rect 15476 12640 15528 12646
rect 14844 9364 14872 9646
rect 15120 9518 15148 12600
rect 15528 12600 15608 12628
rect 15476 12582 15528 12588
rect 15233 12540 15541 12549
rect 15233 12538 15239 12540
rect 15295 12538 15319 12540
rect 15375 12538 15399 12540
rect 15455 12538 15479 12540
rect 15535 12538 15541 12540
rect 15295 12486 15297 12538
rect 15477 12486 15479 12538
rect 15233 12484 15239 12486
rect 15295 12484 15319 12486
rect 15375 12484 15399 12486
rect 15455 12484 15479 12486
rect 15535 12484 15541 12486
rect 15233 12475 15541 12484
rect 15580 12442 15608 12600
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15290 12336 15346 12345
rect 15290 12271 15346 12280
rect 15304 12238 15332 12271
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15672 11898 15700 12786
rect 15764 12782 15792 13262
rect 15856 12850 15884 14962
rect 15948 14498 15976 16594
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 16040 16114 16068 16390
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 16040 14793 16068 14894
rect 16026 14784 16082 14793
rect 16026 14719 16082 14728
rect 15948 14470 16068 14498
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15948 12782 15976 14350
rect 16040 13394 16068 14470
rect 16132 13530 16160 26454
rect 17144 26382 17172 28222
rect 18156 26382 18184 28478
rect 19982 28478 20392 28506
rect 19982 28354 20038 28478
rect 20364 26518 20392 28478
rect 21914 28478 22048 28506
rect 21914 28354 21970 28478
rect 20352 26512 20404 26518
rect 20352 26454 20404 26460
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 16684 23118 16712 26318
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 18512 26308 18564 26314
rect 18512 26250 18564 26256
rect 16764 25696 16816 25702
rect 16764 25638 16816 25644
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16684 22094 16712 23054
rect 16592 22066 16712 22094
rect 16394 19408 16450 19417
rect 16394 19343 16450 19352
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16316 16046 16344 16458
rect 16408 16114 16436 19343
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16224 13530 16252 14282
rect 16408 13938 16436 14894
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16500 13682 16528 17070
rect 16592 13705 16620 22066
rect 16776 21690 16804 25638
rect 16960 24410 16988 26250
rect 18144 25968 18196 25974
rect 18144 25910 18196 25916
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 17132 25696 17184 25702
rect 17132 25638 17184 25644
rect 17052 25265 17080 25638
rect 17038 25256 17094 25265
rect 17038 25191 17094 25200
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16868 21570 16896 23666
rect 16684 21542 16896 21570
rect 16684 20942 16712 21542
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 16684 19446 16712 20878
rect 16672 19440 16724 19446
rect 16672 19382 16724 19388
rect 16684 15094 16712 19382
rect 16868 17202 16896 21422
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16684 14521 16712 15030
rect 16670 14512 16726 14521
rect 16670 14447 16726 14456
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16684 14006 16712 14282
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16684 13734 16712 13806
rect 16672 13728 16724 13734
rect 16316 13654 16528 13682
rect 16578 13696 16634 13705
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16120 13320 16172 13326
rect 16316 13274 16344 13654
rect 16672 13670 16724 13676
rect 16578 13631 16634 13640
rect 16776 13569 16804 16390
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16868 13734 16896 15506
rect 16960 14890 16988 20402
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16762 13560 16818 13569
rect 16762 13495 16818 13504
rect 16580 13456 16632 13462
rect 16578 13424 16580 13433
rect 16632 13424 16634 13433
rect 16578 13359 16634 13368
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16120 13262 16172 13268
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15660 11552 15712 11558
rect 15658 11520 15660 11529
rect 15712 11520 15714 11529
rect 15233 11452 15541 11461
rect 15658 11455 15714 11464
rect 15233 11450 15239 11452
rect 15295 11450 15319 11452
rect 15375 11450 15399 11452
rect 15455 11450 15479 11452
rect 15535 11450 15541 11452
rect 15295 11398 15297 11450
rect 15477 11398 15479 11450
rect 15233 11396 15239 11398
rect 15295 11396 15319 11398
rect 15375 11396 15399 11398
rect 15455 11396 15479 11398
rect 15535 11396 15541 11398
rect 15233 11387 15541 11396
rect 15658 11384 15714 11393
rect 15658 11319 15660 11328
rect 15712 11319 15714 11328
rect 15660 11290 15712 11296
rect 15382 11112 15438 11121
rect 15382 11047 15438 11056
rect 15396 10810 15424 11047
rect 15764 10962 15792 12718
rect 15842 12472 15898 12481
rect 15842 12407 15898 12416
rect 15856 11830 15884 12407
rect 16026 12336 16082 12345
rect 16026 12271 16082 12280
rect 16040 12102 16068 12271
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16040 11218 16068 11698
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15764 10934 15976 10962
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15233 10364 15541 10373
rect 15233 10362 15239 10364
rect 15295 10362 15319 10364
rect 15375 10362 15399 10364
rect 15455 10362 15479 10364
rect 15535 10362 15541 10364
rect 15295 10310 15297 10362
rect 15477 10310 15479 10362
rect 15233 10308 15239 10310
rect 15295 10308 15319 10310
rect 15375 10308 15399 10310
rect 15455 10308 15479 10310
rect 15535 10308 15541 10310
rect 15233 10299 15541 10308
rect 15580 9636 15608 10746
rect 15658 10432 15714 10441
rect 15658 10367 15714 10376
rect 15672 9994 15700 10367
rect 15842 10296 15898 10305
rect 15842 10231 15898 10240
rect 15856 10033 15884 10231
rect 15842 10024 15898 10033
rect 15660 9988 15712 9994
rect 15842 9959 15898 9968
rect 15660 9930 15712 9936
rect 15396 9608 15608 9636
rect 15292 9580 15344 9586
rect 15396 9568 15424 9608
rect 15344 9540 15424 9568
rect 15292 9522 15344 9528
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15488 9450 15516 9608
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 14844 9336 15056 9364
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14832 9104 14884 9110
rect 14738 9072 14794 9081
rect 14884 9064 14964 9092
rect 14832 9046 14884 9052
rect 14738 9007 14794 9016
rect 14752 8838 14780 9007
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14844 8498 14872 8910
rect 14936 8634 14964 9064
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14660 8266 14872 8294
rect 14384 8214 14596 8242
rect 14370 8120 14426 8129
rect 14370 8055 14372 8064
rect 14424 8055 14426 8064
rect 14372 8026 14424 8032
rect 14568 8022 14596 8214
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14292 7206 14320 7686
rect 14476 7478 14504 7686
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 14292 5794 14320 6870
rect 14568 6497 14596 7822
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14752 7002 14780 7414
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14554 6488 14610 6497
rect 14554 6423 14610 6432
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14476 5914 14504 6190
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14568 5914 14596 6122
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14844 5846 14872 8266
rect 14936 7177 14964 8570
rect 15028 7886 15056 9336
rect 15233 9276 15541 9285
rect 15233 9274 15239 9276
rect 15295 9274 15319 9276
rect 15375 9274 15399 9276
rect 15455 9274 15479 9276
rect 15535 9274 15541 9276
rect 15295 9222 15297 9274
rect 15477 9222 15479 9274
rect 15233 9220 15239 9222
rect 15295 9220 15319 9222
rect 15375 9220 15399 9222
rect 15455 9220 15479 9222
rect 15535 9220 15541 9222
rect 15233 9211 15541 9220
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15106 9072 15162 9081
rect 15106 9007 15108 9016
rect 15160 9007 15162 9016
rect 15382 9072 15438 9081
rect 15382 9007 15438 9016
rect 15476 9036 15528 9042
rect 15108 8978 15160 8984
rect 15396 8906 15424 9007
rect 15476 8978 15528 8984
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15304 8276 15332 8774
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15396 8430 15424 8570
rect 15488 8480 15516 8978
rect 15580 8548 15608 9114
rect 15844 9036 15896 9042
rect 15948 9024 15976 10934
rect 16026 10840 16082 10849
rect 16026 10775 16082 10784
rect 16040 9926 16068 10775
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 16040 9625 16068 9862
rect 16132 9722 16160 13262
rect 16224 13246 16344 13274
rect 16224 12170 16252 13246
rect 16316 13110 16620 13138
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 16316 11778 16344 13110
rect 16394 13016 16450 13025
rect 16394 12951 16396 12960
rect 16448 12951 16450 12960
rect 16488 12980 16540 12986
rect 16396 12922 16448 12928
rect 16488 12922 16540 12928
rect 16500 12594 16528 12922
rect 16592 12646 16620 13110
rect 16684 13002 16712 13330
rect 16776 13326 16804 13495
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16764 13184 16816 13190
rect 16762 13152 16764 13161
rect 16816 13152 16818 13161
rect 16762 13087 16818 13096
rect 16684 12986 16804 13002
rect 16684 12980 16816 12986
rect 16684 12974 16764 12980
rect 16764 12922 16816 12928
rect 16408 12566 16528 12594
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16408 12442 16436 12566
rect 16396 12436 16448 12442
rect 16776 12434 16804 12922
rect 16396 12378 16448 12384
rect 16684 12406 16804 12434
rect 16868 12424 16896 13330
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16960 12646 16988 13194
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16488 12300 16540 12306
rect 16684 12288 16712 12406
rect 16868 12396 16988 12424
rect 16540 12260 16712 12288
rect 16764 12300 16816 12306
rect 16488 12242 16540 12248
rect 16764 12242 16816 12248
rect 16776 12102 16804 12242
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16776 11812 16804 12038
rect 16856 11892 16908 11898
rect 16960 11880 16988 12396
rect 16908 11852 16988 11880
rect 16856 11834 16908 11840
rect 16500 11784 16804 11812
rect 16316 11750 16436 11778
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16224 11082 16252 11630
rect 16316 11354 16344 11630
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16210 10976 16266 10985
rect 16210 10911 16266 10920
rect 16224 10577 16252 10911
rect 16210 10568 16266 10577
rect 16210 10503 16266 10512
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16224 9654 16252 9930
rect 16212 9648 16264 9654
rect 16026 9616 16082 9625
rect 16212 9590 16264 9596
rect 16316 9586 16344 9998
rect 16026 9551 16082 9560
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16026 9208 16082 9217
rect 16026 9143 16082 9152
rect 15896 8996 15976 9024
rect 15844 8978 15896 8984
rect 15934 8936 15990 8945
rect 15752 8900 15804 8906
rect 15934 8871 15990 8880
rect 15752 8842 15804 8848
rect 15764 8634 15792 8842
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15580 8520 15700 8548
rect 15488 8452 15608 8480
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15120 8248 15332 8276
rect 15120 8129 15148 8248
rect 15233 8188 15541 8197
rect 15233 8186 15239 8188
rect 15295 8186 15319 8188
rect 15375 8186 15399 8188
rect 15455 8186 15479 8188
rect 15535 8186 15541 8188
rect 15295 8134 15297 8186
rect 15477 8134 15479 8186
rect 15233 8132 15239 8134
rect 15295 8132 15319 8134
rect 15375 8132 15399 8134
rect 15455 8132 15479 8134
rect 15535 8132 15541 8134
rect 15106 8120 15162 8129
rect 15233 8123 15541 8132
rect 15106 8055 15162 8064
rect 15580 7954 15608 8452
rect 15200 7948 15252 7954
rect 15120 7908 15200 7936
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15028 7546 15056 7822
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14922 7168 14978 7177
rect 14922 7103 14978 7112
rect 15028 6798 15056 7482
rect 15120 7002 15148 7908
rect 15200 7890 15252 7896
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15233 7100 15541 7109
rect 15233 7098 15239 7100
rect 15295 7098 15319 7100
rect 15375 7098 15399 7100
rect 15455 7098 15479 7100
rect 15535 7098 15541 7100
rect 15295 7046 15297 7098
rect 15477 7046 15479 7098
rect 15233 7044 15239 7046
rect 15295 7044 15319 7046
rect 15375 7044 15399 7046
rect 15455 7044 15479 7046
rect 15535 7044 15541 7046
rect 15233 7035 15541 7044
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15120 6390 15148 6938
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15396 6730 15424 6870
rect 15672 6780 15700 8520
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15764 8362 15792 8434
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15764 7818 15792 7890
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 15750 7168 15806 7177
rect 15750 7103 15806 7112
rect 15764 6934 15792 7103
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15672 6752 15792 6780
rect 15856 6769 15884 7958
rect 15948 7002 15976 8871
rect 16040 8362 16068 9143
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 15488 6338 15516 6666
rect 15488 6310 15700 6338
rect 15233 6012 15541 6021
rect 15233 6010 15239 6012
rect 15295 6010 15319 6012
rect 15375 6010 15399 6012
rect 15455 6010 15479 6012
rect 15535 6010 15541 6012
rect 15295 5958 15297 6010
rect 15477 5958 15479 6010
rect 15233 5956 15239 5958
rect 15295 5956 15319 5958
rect 15375 5956 15399 5958
rect 15455 5956 15479 5958
rect 15535 5956 15541 5958
rect 14922 5944 14978 5953
rect 15233 5947 15541 5956
rect 14922 5879 14978 5888
rect 14832 5840 14884 5846
rect 14292 5766 14504 5794
rect 14832 5782 14884 5788
rect 14200 5664 14320 5692
rect 14096 5646 14148 5652
rect 14292 5545 14320 5664
rect 14278 5536 14334 5545
rect 14278 5471 14334 5480
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 13832 4678 14044 4706
rect 13832 3534 13860 4678
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 13924 4282 13952 4558
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13924 3233 13952 3946
rect 13910 3224 13966 3233
rect 13910 3159 13966 3168
rect 14016 2854 14044 4218
rect 14108 3942 14136 5170
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14200 4078 14228 4694
rect 14292 4486 14320 5471
rect 14370 4992 14426 5001
rect 14370 4927 14426 4936
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14108 3534 14136 3878
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14188 3120 14240 3126
rect 14094 3088 14150 3097
rect 14292 3108 14320 4082
rect 14384 3126 14412 4927
rect 14476 4622 14504 5766
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14738 5672 14794 5681
rect 14568 4690 14596 5646
rect 14738 5607 14794 5616
rect 14752 5574 14780 5607
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14844 5352 14872 5782
rect 14936 5778 14964 5879
rect 15198 5808 15254 5817
rect 14924 5772 14976 5778
rect 15198 5743 15254 5752
rect 14924 5714 14976 5720
rect 14752 5324 14872 5352
rect 15016 5364 15068 5370
rect 14752 4758 14780 5324
rect 15016 5306 15068 5312
rect 14832 5160 14884 5166
rect 14830 5128 14832 5137
rect 15028 5137 15056 5306
rect 14884 5128 14886 5137
rect 14830 5063 14886 5072
rect 15014 5128 15070 5137
rect 15212 5114 15240 5743
rect 15672 5710 15700 6310
rect 15764 6089 15792 6752
rect 15842 6760 15898 6769
rect 15842 6695 15898 6704
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 15750 6080 15806 6089
rect 15750 6015 15806 6024
rect 15750 5944 15806 5953
rect 15750 5879 15752 5888
rect 15804 5879 15806 5888
rect 15752 5850 15804 5856
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15488 5574 15516 5646
rect 15476 5568 15528 5574
rect 15382 5536 15438 5545
rect 15476 5510 15528 5516
rect 15566 5536 15622 5545
rect 15382 5471 15438 5480
rect 15566 5471 15622 5480
rect 15292 5296 15344 5302
rect 15290 5264 15292 5273
rect 15344 5264 15346 5273
rect 15290 5199 15346 5208
rect 15396 5166 15424 5471
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15488 5273 15516 5306
rect 15474 5264 15530 5273
rect 15474 5199 15530 5208
rect 15014 5063 15070 5072
rect 15120 5086 15240 5114
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14936 4690 14964 4966
rect 15120 4706 15148 5086
rect 15233 4924 15541 4933
rect 15233 4922 15239 4924
rect 15295 4922 15319 4924
rect 15375 4922 15399 4924
rect 15455 4922 15479 4924
rect 15535 4922 15541 4924
rect 15295 4870 15297 4922
rect 15477 4870 15479 4922
rect 15233 4868 15239 4870
rect 15295 4868 15319 4870
rect 15375 4868 15399 4870
rect 15455 4868 15479 4870
rect 15535 4868 15541 4870
rect 15233 4859 15541 4868
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14924 4684 14976 4690
rect 15120 4678 15240 4706
rect 14924 4626 14976 4632
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14554 4584 14610 4593
rect 14554 4519 14556 4528
rect 14608 4519 14610 4528
rect 14556 4490 14608 4496
rect 14832 4208 14884 4214
rect 14936 4162 14964 4626
rect 15212 4214 15240 4678
rect 15580 4554 15608 5471
rect 15672 5370 15700 5646
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15672 4690 15700 5306
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 14884 4156 14964 4162
rect 14832 4150 14964 4156
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 14844 4134 14964 4150
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14660 3670 14688 4014
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14936 3602 14964 4134
rect 15488 3924 15516 4490
rect 15566 4312 15622 4321
rect 15566 4247 15622 4256
rect 15580 4078 15608 4247
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15752 3936 15804 3942
rect 15488 3896 15752 3924
rect 15752 3878 15804 3884
rect 15233 3836 15541 3845
rect 15233 3834 15239 3836
rect 15295 3834 15319 3836
rect 15375 3834 15399 3836
rect 15455 3834 15479 3836
rect 15535 3834 15541 3836
rect 15295 3782 15297 3834
rect 15477 3782 15479 3834
rect 15233 3780 15239 3782
rect 15295 3780 15319 3782
rect 15375 3780 15399 3782
rect 15455 3780 15479 3782
rect 15535 3780 15541 3782
rect 15233 3771 15541 3780
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15488 3194 15516 3402
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 14240 3080 14320 3108
rect 14188 3062 14240 3068
rect 14094 3023 14150 3032
rect 14108 2854 14136 3023
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 13740 2746 13952 2774
rect 13818 2272 13874 2281
rect 13818 2207 13874 2216
rect 13634 2136 13690 2145
rect 13832 2106 13860 2207
rect 13634 2071 13690 2080
rect 13820 2100 13872 2106
rect 13820 2042 13872 2048
rect 13544 1896 13596 1902
rect 13544 1838 13596 1844
rect 13266 1728 13322 1737
rect 13266 1663 13322 1672
rect 10232 128 10284 134
rect 10232 70 10284 76
rect 10322 0 10378 800
rect 12254 0 12310 800
rect 13924 762 13952 2746
rect 14292 2514 14320 3080
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 15233 2748 15541 2757
rect 15233 2746 15239 2748
rect 15295 2746 15319 2748
rect 15375 2746 15399 2748
rect 15455 2746 15479 2748
rect 15535 2746 15541 2748
rect 15295 2694 15297 2746
rect 15477 2694 15479 2746
rect 15233 2692 15239 2694
rect 15295 2692 15319 2694
rect 15375 2692 15399 2694
rect 15455 2692 15479 2694
rect 15535 2692 15541 2694
rect 15233 2683 15541 2692
rect 15856 2650 15884 6326
rect 15948 5778 15976 6598
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16040 5642 16068 6122
rect 16224 5953 16252 9386
rect 16408 9058 16436 11750
rect 16500 10606 16528 11784
rect 17052 11762 17080 24550
rect 17144 17270 17172 25638
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17316 24880 17368 24886
rect 17316 24822 17368 24828
rect 17224 24268 17276 24274
rect 17224 24210 17276 24216
rect 17236 21622 17264 24210
rect 17328 23730 17356 24822
rect 17684 24744 17736 24750
rect 17684 24686 17736 24692
rect 17408 24676 17460 24682
rect 17408 24618 17460 24624
rect 17420 23730 17448 24618
rect 17696 23730 17724 24686
rect 17880 24410 17908 25298
rect 18156 25294 18184 25910
rect 18524 25906 18552 26250
rect 19994 26140 20302 26149
rect 19994 26138 20000 26140
rect 20056 26138 20080 26140
rect 20136 26138 20160 26140
rect 20216 26138 20240 26140
rect 20296 26138 20302 26140
rect 20056 26086 20058 26138
rect 20238 26086 20240 26138
rect 19994 26084 20000 26086
rect 20056 26084 20080 26086
rect 20136 26084 20160 26086
rect 20216 26084 20240 26086
rect 20296 26084 20302 26086
rect 19994 26075 20302 26084
rect 18880 26036 18932 26042
rect 18880 25978 18932 25984
rect 18512 25900 18564 25906
rect 18512 25842 18564 25848
rect 18236 25832 18288 25838
rect 18236 25774 18288 25780
rect 18248 25362 18276 25774
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18156 24818 18184 25094
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 18156 24274 18184 24754
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17420 20398 17448 23666
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17696 19854 17724 23666
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17880 22094 17908 23462
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 17972 22098 18000 22646
rect 17788 22066 17908 22094
rect 17960 22092 18012 22098
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17788 19786 17816 22066
rect 17960 22034 18012 22040
rect 17776 19780 17828 19786
rect 17776 19722 17828 19728
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17236 16794 17264 19314
rect 17512 18358 17540 19654
rect 17788 18698 17816 19722
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18248 19334 18276 25298
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17500 18352 17552 18358
rect 17406 18320 17462 18329
rect 17500 18294 17552 18300
rect 17880 18290 17908 18634
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 17406 18255 17462 18264
rect 17592 18284 17644 18290
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17236 16590 17264 16730
rect 17328 16590 17356 17546
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17236 14958 17264 16526
rect 17314 16008 17370 16017
rect 17314 15943 17370 15952
rect 17328 15337 17356 15943
rect 17314 15328 17370 15337
rect 17314 15263 17370 15272
rect 17420 15144 17448 18255
rect 17592 18226 17644 18232
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17328 15116 17448 15144
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16578 11112 16634 11121
rect 16578 11047 16634 11056
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16500 9722 16528 10134
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16486 9616 16542 9625
rect 16486 9551 16488 9560
rect 16540 9551 16542 9560
rect 16488 9522 16540 9528
rect 16316 9030 16436 9058
rect 16316 8090 16344 9030
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16408 7206 16436 8366
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16394 7032 16450 7041
rect 16394 6967 16450 6976
rect 16408 6866 16436 6967
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16500 6497 16528 9522
rect 16592 7818 16620 11047
rect 16684 10742 16712 11494
rect 17144 11354 17172 13466
rect 17236 12374 17264 13738
rect 17328 12374 17356 15116
rect 17512 15094 17540 17478
rect 17500 15088 17552 15094
rect 17406 15056 17462 15065
rect 17500 15030 17552 15036
rect 17406 14991 17462 15000
rect 17420 13870 17448 14991
rect 17500 14952 17552 14958
rect 17498 14920 17500 14929
rect 17552 14920 17554 14929
rect 17498 14855 17554 14864
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17420 12306 17448 13466
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17512 12186 17540 14554
rect 17604 14346 17632 18226
rect 17880 18193 17908 18226
rect 17866 18184 17922 18193
rect 17866 18119 17922 18128
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17880 15978 17908 18022
rect 17972 16794 18000 18362
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17972 15502 18000 16390
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17420 12158 17540 12186
rect 17420 11937 17448 12158
rect 17498 12064 17554 12073
rect 17498 11999 17554 12008
rect 17406 11928 17462 11937
rect 17406 11863 17462 11872
rect 17512 11830 17540 11999
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17408 11756 17460 11762
rect 17328 11716 17408 11744
rect 17328 11354 17356 11716
rect 17408 11698 17460 11704
rect 17498 11520 17554 11529
rect 17498 11455 17554 11464
rect 17512 11354 17540 11455
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 16946 11112 17002 11121
rect 16946 11047 17002 11056
rect 16764 11008 16816 11014
rect 16960 10996 16988 11047
rect 17132 11008 17184 11014
rect 16764 10950 16816 10956
rect 16868 10968 17132 10996
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 16776 10198 16804 10950
rect 16868 10418 16896 10968
rect 17132 10950 17184 10956
rect 17328 10606 17356 11290
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17420 10606 17448 11154
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17132 10464 17184 10470
rect 16868 10390 16988 10418
rect 17132 10406 17184 10412
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16776 9586 16804 9998
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16776 8498 16804 9522
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16684 8294 16712 8434
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16776 8106 16804 8434
rect 16684 8078 16804 8106
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16684 6934 16712 8078
rect 16762 7984 16818 7993
rect 16868 7954 16896 9658
rect 16762 7919 16764 7928
rect 16816 7919 16818 7928
rect 16856 7948 16908 7954
rect 16764 7890 16816 7896
rect 16856 7890 16908 7896
rect 16776 7478 16804 7890
rect 16960 7585 16988 10390
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 17052 8566 17080 9590
rect 17144 8566 17172 10406
rect 17224 9920 17276 9926
rect 17222 9888 17224 9897
rect 17276 9888 17278 9897
rect 17222 9823 17278 9832
rect 17328 9674 17356 10542
rect 17512 10538 17540 10678
rect 17500 10532 17552 10538
rect 17500 10474 17552 10480
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17236 9646 17356 9674
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17236 8412 17264 9646
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 8809 17356 9318
rect 17314 8800 17370 8809
rect 17314 8735 17370 8744
rect 17038 8392 17094 8401
rect 17038 8327 17094 8336
rect 17144 8384 17264 8412
rect 16946 7576 17002 7585
rect 17052 7546 17080 8327
rect 16946 7511 17002 7520
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16948 7472 17000 7478
rect 17144 7426 17172 8384
rect 17222 8120 17278 8129
rect 17222 8055 17278 8064
rect 17236 7449 17264 8055
rect 17314 7576 17370 7585
rect 17314 7511 17370 7520
rect 16948 7414 17000 7420
rect 16672 6928 16724 6934
rect 16672 6870 16724 6876
rect 16960 6730 16988 7414
rect 17052 7398 17172 7426
rect 17222 7440 17278 7449
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16486 6488 16542 6497
rect 16486 6423 16542 6432
rect 16578 6352 16634 6361
rect 16578 6287 16634 6296
rect 16592 6118 16620 6287
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16210 5944 16266 5953
rect 16210 5879 16266 5888
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 16670 5536 16726 5545
rect 16670 5471 16726 5480
rect 16118 5264 16174 5273
rect 16118 5199 16174 5208
rect 16132 5098 16160 5199
rect 16120 5092 16172 5098
rect 16120 5034 16172 5040
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16316 4729 16344 4966
rect 16580 4752 16632 4758
rect 16302 4720 16358 4729
rect 16580 4694 16632 4700
rect 16302 4655 16358 4664
rect 16302 4176 16358 4185
rect 16302 4111 16304 4120
rect 16356 4111 16358 4120
rect 16304 4082 16356 4088
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15198 2544 15254 2553
rect 14280 2508 14332 2514
rect 15198 2479 15254 2488
rect 14280 2450 14332 2456
rect 15212 2378 15240 2479
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 14568 1698 14596 2314
rect 14556 1692 14608 1698
rect 14556 1634 14608 1640
rect 15948 950 15976 2994
rect 16316 2774 16344 3674
rect 16592 3602 16620 4694
rect 16684 4622 16712 5471
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16224 2746 16344 2774
rect 16224 1562 16252 2746
rect 16500 1970 16528 3402
rect 16868 3058 16896 3538
rect 16960 3398 16988 4558
rect 17052 4146 17080 7398
rect 17328 7410 17356 7511
rect 17222 7375 17278 7384
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17420 7290 17448 10066
rect 17604 9602 17632 13942
rect 17696 13734 17724 15302
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17880 14618 17908 14826
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 14385 17908 14418
rect 17866 14376 17922 14385
rect 17866 14311 17922 14320
rect 17972 14260 18000 15302
rect 18064 15162 18092 17682
rect 18156 17270 18184 19314
rect 18248 19306 18368 19334
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18156 15042 18184 16730
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 17880 14232 18000 14260
rect 18064 15014 18184 15042
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17788 13530 17816 13670
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17696 12374 17724 13194
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17788 12442 17816 12582
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17684 12368 17736 12374
rect 17684 12310 17736 12316
rect 17774 12336 17830 12345
rect 17774 12271 17830 12280
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11937 17724 12174
rect 17682 11928 17738 11937
rect 17682 11863 17738 11872
rect 17788 11778 17816 12271
rect 17880 12170 17908 14232
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17866 12064 17922 12073
rect 17866 11999 17922 12008
rect 17696 11750 17816 11778
rect 17880 11762 17908 11999
rect 17972 11898 18000 12310
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17868 11756 17920 11762
rect 17696 10130 17724 11750
rect 17868 11698 17920 11704
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17774 11656 17830 11665
rect 17774 11591 17830 11600
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17788 9654 17816 11591
rect 17880 11393 17908 11698
rect 17866 11384 17922 11393
rect 17866 11319 17922 11328
rect 17972 11150 18000 11698
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17776 9648 17828 9654
rect 17604 9574 17724 9602
rect 17776 9590 17828 9596
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17604 8974 17632 9454
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17512 8673 17540 8842
rect 17498 8664 17554 8673
rect 17498 8599 17554 8608
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17512 7818 17540 8230
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17498 7712 17554 7721
rect 17498 7647 17554 7656
rect 17328 7262 17448 7290
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17144 7002 17172 7142
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17236 5556 17264 6394
rect 17328 5710 17356 7262
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17316 5568 17368 5574
rect 17236 5528 17316 5556
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17144 4826 17172 5238
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17236 4146 17264 5528
rect 17316 5510 17368 5516
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 17144 3602 17172 3946
rect 17328 3942 17356 4082
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17038 3496 17094 3505
rect 17420 3466 17448 7142
rect 17512 6730 17540 7647
rect 17604 7041 17632 8502
rect 17590 7032 17646 7041
rect 17590 6967 17646 6976
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17498 6488 17554 6497
rect 17498 6423 17554 6432
rect 17512 6322 17540 6423
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17038 3431 17094 3440
rect 17408 3460 17460 3466
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16488 1964 16540 1970
rect 16488 1906 16540 1912
rect 16776 1834 16804 2926
rect 16868 2514 16896 2994
rect 17052 2825 17080 3431
rect 17408 3402 17460 3408
rect 17038 2816 17094 2825
rect 17038 2751 17094 2760
rect 17130 2680 17186 2689
rect 17130 2615 17186 2624
rect 17144 2514 17172 2615
rect 17512 2514 17540 6258
rect 17590 6080 17646 6089
rect 17590 6015 17646 6024
rect 17604 5302 17632 6015
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17604 4214 17632 4762
rect 17696 4690 17724 9574
rect 17788 9489 17816 9590
rect 17880 9518 17908 10542
rect 17972 9722 18000 11086
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17868 9512 17920 9518
rect 17774 9480 17830 9489
rect 17868 9454 17920 9460
rect 17774 9415 17830 9424
rect 17776 8084 17828 8090
rect 17960 8084 18012 8090
rect 17828 8044 17908 8072
rect 17776 8026 17828 8032
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17788 5914 17816 7822
rect 17880 7206 17908 8044
rect 17960 8026 18012 8032
rect 17972 7886 18000 8026
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7342 18000 7686
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17958 6624 18014 6633
rect 17958 6559 18014 6568
rect 17972 6458 18000 6559
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17880 5370 17908 6190
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17972 5370 18000 5510
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17880 4146 17908 5306
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17958 4040 18014 4049
rect 17788 3602 17816 4014
rect 17958 3975 18014 3984
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17972 3466 18000 3975
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17868 2644 17920 2650
rect 18064 2632 18092 15014
rect 18248 13938 18276 15098
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18248 13258 18276 13738
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18156 8090 18184 13194
rect 18340 12730 18368 19306
rect 18432 15042 18460 22578
rect 18524 15162 18552 25842
rect 18604 25220 18656 25226
rect 18604 25162 18656 25168
rect 18616 24954 18644 25162
rect 18604 24948 18656 24954
rect 18604 24890 18656 24896
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18616 23050 18644 24210
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18616 22166 18644 22986
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 18708 22030 18736 22510
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18708 20777 18736 21830
rect 18694 20768 18750 20777
rect 18694 20703 18750 20712
rect 18800 20262 18828 22714
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18708 16833 18736 19790
rect 18800 19378 18828 20198
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18892 18442 18920 25978
rect 19994 25052 20302 25061
rect 19994 25050 20000 25052
rect 20056 25050 20080 25052
rect 20136 25050 20160 25052
rect 20216 25050 20240 25052
rect 20296 25050 20302 25052
rect 20056 24998 20058 25050
rect 20238 24998 20240 25050
rect 19994 24996 20000 24998
rect 20056 24996 20080 24998
rect 20136 24996 20160 24998
rect 20216 24996 20240 24998
rect 20296 24996 20302 24998
rect 19994 24987 20302 24996
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 19076 22778 19104 24278
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19156 23248 19208 23254
rect 19156 23190 19208 23196
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 18984 21486 19012 21898
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 19168 21049 19196 23190
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19260 21962 19288 23122
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 19248 21956 19300 21962
rect 19248 21898 19300 21904
rect 19154 21040 19210 21049
rect 19154 20975 19210 20984
rect 19352 19961 19380 22442
rect 19720 22094 19748 24006
rect 19994 23964 20302 23973
rect 19994 23962 20000 23964
rect 20056 23962 20080 23964
rect 20136 23962 20160 23964
rect 20216 23962 20240 23964
rect 20296 23962 20302 23964
rect 20056 23910 20058 23962
rect 20238 23910 20240 23962
rect 19994 23908 20000 23910
rect 20056 23908 20080 23910
rect 20136 23908 20160 23910
rect 20216 23908 20240 23910
rect 20296 23908 20302 23910
rect 19994 23899 20302 23908
rect 19994 22876 20302 22885
rect 19994 22874 20000 22876
rect 20056 22874 20080 22876
rect 20136 22874 20160 22876
rect 20216 22874 20240 22876
rect 20296 22874 20302 22876
rect 20056 22822 20058 22874
rect 20238 22822 20240 22874
rect 19994 22820 20000 22822
rect 20056 22820 20080 22822
rect 20136 22820 20160 22822
rect 20216 22820 20240 22822
rect 20296 22820 20302 22822
rect 19994 22811 20302 22820
rect 19628 22066 19748 22094
rect 19338 19952 19394 19961
rect 19338 19887 19394 19896
rect 19294 19848 19346 19854
rect 19346 19808 19564 19836
rect 19294 19790 19346 19796
rect 19536 19718 19564 19808
rect 19248 19712 19300 19718
rect 19524 19712 19576 19718
rect 19248 19654 19300 19660
rect 19338 19680 19394 19689
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18800 18414 18920 18442
rect 18800 17134 18828 18414
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18694 16824 18750 16833
rect 18694 16759 18750 16768
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18432 15014 18552 15042
rect 18420 14816 18472 14822
rect 18524 14793 18552 15014
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18420 14758 18472 14764
rect 18510 14784 18566 14793
rect 18432 13530 18460 14758
rect 18510 14719 18566 14728
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18248 12702 18368 12730
rect 18248 11762 18276 12702
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18248 11286 18276 11494
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 8974 18276 9318
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18340 7698 18368 12582
rect 18432 12186 18460 13194
rect 18524 13025 18552 14282
rect 18616 14113 18644 14894
rect 18602 14104 18658 14113
rect 18602 14039 18658 14048
rect 18510 13016 18566 13025
rect 18510 12951 18566 12960
rect 18616 12646 18644 14039
rect 18708 13326 18736 16759
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18800 13802 18828 14486
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18786 13560 18842 13569
rect 18786 13495 18788 13504
rect 18840 13495 18842 13504
rect 18788 13466 18840 13472
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18892 13240 18920 18226
rect 18800 13212 18920 13240
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18708 12306 18736 12922
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18432 12158 18552 12186
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11558 18460 12038
rect 18524 11830 18552 12158
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18248 7670 18368 7698
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 18156 5846 18184 7210
rect 18248 6866 18276 7670
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18340 7002 18368 7482
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 18340 5710 18368 6938
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18340 4321 18368 4626
rect 18326 4312 18382 4321
rect 18326 4247 18382 4256
rect 18234 4040 18290 4049
rect 18234 3975 18290 3984
rect 18248 3058 18276 3975
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18144 2644 18196 2650
rect 18064 2604 18144 2632
rect 17868 2586 17920 2592
rect 18144 2586 18196 2592
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17236 2310 17264 2450
rect 17880 2310 17908 2586
rect 18432 2378 18460 11290
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18524 10266 18552 11018
rect 18616 10985 18644 11698
rect 18602 10976 18658 10985
rect 18602 10911 18658 10920
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18616 8906 18644 10746
rect 18708 9761 18736 11834
rect 18800 10470 18828 13212
rect 18984 13172 19012 19314
rect 19156 15428 19208 15434
rect 19156 15370 19208 15376
rect 18892 13144 19012 13172
rect 18892 12986 18920 13144
rect 19062 13016 19118 13025
rect 18880 12980 18932 12986
rect 19062 12951 19118 12960
rect 18880 12922 18932 12928
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18984 11898 19012 12854
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18694 9752 18750 9761
rect 18694 9687 18750 9696
rect 18708 8974 18736 9687
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18524 6390 18552 8298
rect 18708 7886 18736 8774
rect 18800 8480 18828 10406
rect 19076 9674 19104 12951
rect 19168 12186 19196 15370
rect 19260 15042 19288 19654
rect 19524 19654 19576 19660
rect 19338 19615 19394 19624
rect 19352 17377 19380 19615
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19444 18426 19472 19314
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19536 18358 19564 18634
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19338 17368 19394 17377
rect 19338 17303 19394 17312
rect 19536 16969 19564 18294
rect 19522 16960 19578 16969
rect 19522 16895 19578 16904
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 15094 19472 15302
rect 19432 15088 19484 15094
rect 19260 15014 19380 15042
rect 19432 15030 19484 15036
rect 19352 12306 19380 15014
rect 19432 14952 19484 14958
rect 19430 14920 19432 14929
rect 19484 14920 19486 14929
rect 19430 14855 19486 14864
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19444 13326 19472 13738
rect 19536 13326 19564 16895
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19168 12158 19380 12186
rect 19352 10062 19380 12158
rect 19444 11014 19472 13262
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 18984 9646 19104 9674
rect 18880 8492 18932 8498
rect 18800 8452 18880 8480
rect 18880 8434 18932 8440
rect 18984 8242 19012 9646
rect 19536 9625 19564 11698
rect 19628 11354 19656 22066
rect 19994 21788 20302 21797
rect 19994 21786 20000 21788
rect 20056 21786 20080 21788
rect 20136 21786 20160 21788
rect 20216 21786 20240 21788
rect 20296 21786 20302 21788
rect 20056 21734 20058 21786
rect 20238 21734 20240 21786
rect 19994 21732 20000 21734
rect 20056 21732 20080 21734
rect 20136 21732 20160 21734
rect 20216 21732 20240 21734
rect 20296 21732 20302 21734
rect 19994 21723 20302 21732
rect 19708 21412 19760 21418
rect 19708 21354 19760 21360
rect 19720 19334 19748 21354
rect 19994 20700 20302 20709
rect 19994 20698 20000 20700
rect 20056 20698 20080 20700
rect 20136 20698 20160 20700
rect 20216 20698 20240 20700
rect 20296 20698 20302 20700
rect 20056 20646 20058 20698
rect 20238 20646 20240 20698
rect 19994 20644 20000 20646
rect 20056 20644 20080 20646
rect 20136 20644 20160 20646
rect 20216 20644 20240 20646
rect 20296 20644 20302 20646
rect 19994 20635 20302 20644
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 19812 19786 19840 20538
rect 20352 19984 20404 19990
rect 20352 19926 20404 19932
rect 19890 19816 19946 19825
rect 19800 19780 19852 19786
rect 19890 19751 19946 19760
rect 19800 19722 19852 19728
rect 19812 19446 19840 19722
rect 19904 19446 19932 19751
rect 19994 19612 20302 19621
rect 19994 19610 20000 19612
rect 20056 19610 20080 19612
rect 20136 19610 20160 19612
rect 20216 19610 20240 19612
rect 20296 19610 20302 19612
rect 20056 19558 20058 19610
rect 20238 19558 20240 19610
rect 19994 19556 20000 19558
rect 20056 19556 20080 19558
rect 20136 19556 20160 19558
rect 20216 19556 20240 19558
rect 20296 19556 20302 19558
rect 19994 19547 20302 19556
rect 19800 19440 19852 19446
rect 19800 19382 19852 19388
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 19720 19306 19932 19334
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19720 15434 19748 18702
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19812 17338 19840 17478
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19706 15192 19762 15201
rect 19706 15127 19762 15136
rect 19720 14006 19748 15127
rect 19708 14000 19760 14006
rect 19708 13942 19760 13948
rect 19812 13462 19840 17274
rect 19904 15994 19932 19306
rect 19994 18524 20302 18533
rect 19994 18522 20000 18524
rect 20056 18522 20080 18524
rect 20136 18522 20160 18524
rect 20216 18522 20240 18524
rect 20296 18522 20302 18524
rect 20056 18470 20058 18522
rect 20238 18470 20240 18522
rect 19994 18468 20000 18470
rect 20056 18468 20080 18470
rect 20136 18468 20160 18470
rect 20216 18468 20240 18470
rect 20296 18468 20302 18470
rect 19994 18459 20302 18468
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19996 17542 20024 18226
rect 20364 17678 20392 19926
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20456 18086 20484 19382
rect 20548 19378 20576 24210
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20548 18290 20576 19110
rect 20640 18426 20668 26386
rect 22020 26382 22048 28478
rect 23202 28478 23336 28506
rect 23202 28354 23258 28478
rect 23308 26382 23336 28478
rect 25134 28354 25190 29154
rect 27066 28506 27122 29154
rect 27066 28478 27384 28506
rect 27066 28354 27122 28478
rect 23756 26852 23808 26858
rect 23756 26794 23808 26800
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 23572 26308 23624 26314
rect 23572 26250 23624 26256
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20916 23497 20944 25434
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 20902 23488 20958 23497
rect 20902 23423 20958 23432
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21284 20369 21312 20402
rect 21270 20360 21326 20369
rect 21088 20324 21140 20330
rect 21270 20295 21326 20304
rect 21088 20266 21140 20272
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20732 19689 20760 19790
rect 20718 19680 20774 19689
rect 20718 19615 20774 19624
rect 21100 19514 21128 20266
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21192 19990 21220 20198
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20732 18970 20760 19314
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21192 19174 21220 19246
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19994 17436 20302 17445
rect 19994 17434 20000 17436
rect 20056 17434 20080 17436
rect 20136 17434 20160 17436
rect 20216 17434 20240 17436
rect 20296 17434 20302 17436
rect 20056 17382 20058 17434
rect 20238 17382 20240 17434
rect 19994 17380 20000 17382
rect 20056 17380 20080 17382
rect 20136 17380 20160 17382
rect 20216 17380 20240 17382
rect 20296 17380 20302 17382
rect 19994 17371 20302 17380
rect 19994 16348 20302 16357
rect 19994 16346 20000 16348
rect 20056 16346 20080 16348
rect 20136 16346 20160 16348
rect 20216 16346 20240 16348
rect 20296 16346 20302 16348
rect 20056 16294 20058 16346
rect 20238 16294 20240 16346
rect 19994 16292 20000 16294
rect 20056 16292 20080 16294
rect 20136 16292 20160 16294
rect 20216 16292 20240 16294
rect 20296 16292 20302 16294
rect 19994 16283 20302 16292
rect 20074 16144 20130 16153
rect 20364 16114 20392 17614
rect 20442 16144 20498 16153
rect 20074 16079 20130 16088
rect 20352 16108 20404 16114
rect 19904 15966 20024 15994
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19904 14414 19932 15846
rect 19996 15638 20024 15966
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 20088 15434 20116 16079
rect 20442 16079 20498 16088
rect 20352 16050 20404 16056
rect 20364 15502 20392 16050
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 19994 15260 20302 15269
rect 19994 15258 20000 15260
rect 20056 15258 20080 15260
rect 20136 15258 20160 15260
rect 20216 15258 20240 15260
rect 20296 15258 20302 15260
rect 20056 15206 20058 15258
rect 20238 15206 20240 15258
rect 19994 15204 20000 15206
rect 20056 15204 20080 15206
rect 20136 15204 20160 15206
rect 20216 15204 20240 15206
rect 20296 15204 20302 15206
rect 19994 15195 20302 15204
rect 19984 15088 20036 15094
rect 19982 15056 19984 15065
rect 20036 15056 20038 15065
rect 19982 14991 20038 15000
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19994 14172 20302 14181
rect 19994 14170 20000 14172
rect 20056 14170 20080 14172
rect 20136 14170 20160 14172
rect 20216 14170 20240 14172
rect 20296 14170 20302 14172
rect 20056 14118 20058 14170
rect 20238 14118 20240 14170
rect 19994 14116 20000 14118
rect 20056 14116 20080 14118
rect 20136 14116 20160 14118
rect 20216 14116 20240 14118
rect 20296 14116 20302 14118
rect 19994 14107 20302 14116
rect 20364 14056 20392 15438
rect 19904 14028 20392 14056
rect 19800 13456 19852 13462
rect 19706 13424 19762 13433
rect 19800 13398 19852 13404
rect 19706 13359 19762 13368
rect 19720 12374 19748 13359
rect 19904 13274 19932 14028
rect 20456 13938 20484 16079
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 19812 13246 19932 13274
rect 20444 13252 20496 13258
rect 19708 12368 19760 12374
rect 19708 12310 19760 12316
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19720 10554 19748 11630
rect 19812 10674 19840 13246
rect 20444 13194 20496 13200
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19720 10526 19840 10554
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19522 9616 19578 9625
rect 19522 9551 19578 9560
rect 19720 9518 19748 10066
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19062 9344 19118 9353
rect 19062 9279 19118 9288
rect 18892 8214 19012 8242
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18786 7848 18842 7857
rect 18604 7812 18656 7818
rect 18786 7783 18788 7792
rect 18604 7754 18656 7760
rect 18840 7783 18842 7792
rect 18788 7754 18840 7760
rect 18616 7410 18644 7754
rect 18892 7478 18920 8214
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18524 3738 18552 4422
rect 18616 3738 18644 7346
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18708 5778 18736 6802
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18708 2553 18736 5238
rect 18800 4457 18828 6666
rect 18984 6254 19012 8026
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 19076 5574 19104 9279
rect 19522 9208 19578 9217
rect 19522 9143 19578 9152
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8945 19380 8978
rect 19338 8936 19394 8945
rect 19338 8871 19394 8880
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19444 8362 19472 8774
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19352 7410 19380 7822
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19352 6934 19380 7346
rect 19340 6928 19392 6934
rect 19340 6870 19392 6876
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19076 5030 19104 5102
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19352 4570 19380 5646
rect 19444 5114 19472 7958
rect 19536 6882 19564 9143
rect 19720 8974 19748 9454
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19706 8800 19762 8809
rect 19706 8735 19762 8744
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19628 7750 19656 8230
rect 19720 7857 19748 8735
rect 19812 8412 19840 10526
rect 19904 9926 19932 13126
rect 19994 13084 20302 13093
rect 19994 13082 20000 13084
rect 20056 13082 20080 13084
rect 20136 13082 20160 13084
rect 20216 13082 20240 13084
rect 20296 13082 20302 13084
rect 20056 13030 20058 13082
rect 20238 13030 20240 13082
rect 19994 13028 20000 13030
rect 20056 13028 20080 13030
rect 20136 13028 20160 13030
rect 20216 13028 20240 13030
rect 20296 13028 20302 13030
rect 19994 13019 20302 13028
rect 20364 12442 20392 13126
rect 20456 12646 20484 13194
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 19994 11996 20302 12005
rect 19994 11994 20000 11996
rect 20056 11994 20080 11996
rect 20136 11994 20160 11996
rect 20216 11994 20240 11996
rect 20296 11994 20302 11996
rect 20056 11942 20058 11994
rect 20238 11942 20240 11994
rect 19994 11940 20000 11942
rect 20056 11940 20080 11942
rect 20136 11940 20160 11942
rect 20216 11940 20240 11942
rect 20296 11940 20302 11942
rect 19994 11931 20302 11940
rect 20456 11898 20484 12582
rect 20548 12238 20576 17614
rect 20732 16522 20760 18906
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 21100 17814 21128 18634
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 20640 15026 20668 15574
rect 20732 15502 20760 15982
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20628 14884 20680 14890
rect 20628 14826 20680 14832
rect 20640 14482 20668 14826
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20732 14414 20760 15438
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20732 14006 20760 14350
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20640 12186 20668 13806
rect 20732 13394 20760 13942
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20732 12986 20760 13330
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20720 12232 20772 12238
rect 20640 12180 20720 12186
rect 20640 12174 20772 12180
rect 20640 12158 20760 12174
rect 20824 12170 20852 17070
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 21008 16794 21036 16934
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21008 16658 21036 16730
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20904 15428 20956 15434
rect 20904 15370 20956 15376
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 19994 10908 20302 10917
rect 19994 10906 20000 10908
rect 20056 10906 20080 10908
rect 20136 10906 20160 10908
rect 20216 10906 20240 10908
rect 20296 10906 20302 10908
rect 20056 10854 20058 10906
rect 20238 10854 20240 10906
rect 19994 10852 20000 10854
rect 20056 10852 20080 10854
rect 20136 10852 20160 10854
rect 20216 10852 20240 10854
rect 20296 10852 20302 10854
rect 19994 10843 20302 10852
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19994 9820 20302 9829
rect 19994 9818 20000 9820
rect 20056 9818 20080 9820
rect 20136 9818 20160 9820
rect 20216 9818 20240 9820
rect 20296 9818 20302 9820
rect 20056 9766 20058 9818
rect 20238 9766 20240 9818
rect 19994 9764 20000 9766
rect 20056 9764 20080 9766
rect 20136 9764 20160 9766
rect 20216 9764 20240 9766
rect 20296 9764 20302 9766
rect 19994 9755 20302 9764
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 19904 8514 19932 9658
rect 20352 9648 20404 9654
rect 19982 9616 20038 9625
rect 20352 9590 20404 9596
rect 19982 9551 20038 9560
rect 19996 8974 20024 9551
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19994 8732 20302 8741
rect 19994 8730 20000 8732
rect 20056 8730 20080 8732
rect 20136 8730 20160 8732
rect 20216 8730 20240 8732
rect 20296 8730 20302 8732
rect 20056 8678 20058 8730
rect 20238 8678 20240 8730
rect 19994 8676 20000 8678
rect 20056 8676 20080 8678
rect 20136 8676 20160 8678
rect 20216 8676 20240 8678
rect 20296 8676 20302 8678
rect 19994 8667 20302 8676
rect 19904 8486 20024 8514
rect 20364 8498 20392 9590
rect 20456 9586 20484 11698
rect 20548 11150 20576 11834
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20640 10674 20668 12038
rect 20732 11558 20760 12158
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20732 11218 20760 11494
rect 20720 11212 20772 11218
rect 20772 11172 20852 11200
rect 20720 11154 20772 11160
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20628 10532 20680 10538
rect 20628 10474 20680 10480
rect 20640 10130 20668 10474
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20732 10169 20760 10202
rect 20718 10160 20774 10169
rect 20628 10124 20680 10130
rect 20548 10084 20628 10112
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20548 9042 20576 10084
rect 20718 10095 20774 10104
rect 20628 10066 20680 10072
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 19892 8424 19944 8430
rect 19812 8384 19892 8412
rect 19892 8366 19944 8372
rect 19800 8288 19852 8294
rect 19800 8230 19852 8236
rect 19706 7848 19762 7857
rect 19706 7783 19762 7792
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19812 7041 19840 8230
rect 19996 7732 20024 8486
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 20272 7750 20300 8298
rect 19904 7704 20024 7732
rect 20260 7744 20312 7750
rect 19798 7032 19854 7041
rect 19798 6967 19854 6976
rect 19536 6854 19656 6882
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19536 5522 19564 6734
rect 19628 5914 19656 6854
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19720 6254 19748 6666
rect 19904 6440 19932 7704
rect 20260 7686 20312 7692
rect 19994 7644 20302 7653
rect 19994 7642 20000 7644
rect 20056 7642 20080 7644
rect 20136 7642 20160 7644
rect 20216 7642 20240 7644
rect 20296 7642 20302 7644
rect 20056 7590 20058 7642
rect 20238 7590 20240 7642
rect 19994 7588 20000 7590
rect 20056 7588 20080 7590
rect 20136 7588 20160 7590
rect 20216 7588 20240 7590
rect 20296 7588 20302 7590
rect 19994 7579 20302 7588
rect 19994 6556 20302 6565
rect 19994 6554 20000 6556
rect 20056 6554 20080 6556
rect 20136 6554 20160 6556
rect 20216 6554 20240 6556
rect 20296 6554 20302 6556
rect 20056 6502 20058 6554
rect 20238 6502 20240 6554
rect 19994 6500 20000 6502
rect 20056 6500 20080 6502
rect 20136 6500 20160 6502
rect 20216 6500 20240 6502
rect 20296 6500 20302 6502
rect 19994 6491 20302 6500
rect 19904 6412 20024 6440
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19720 5846 19748 6190
rect 19708 5840 19760 5846
rect 19614 5808 19670 5817
rect 19708 5782 19760 5788
rect 19614 5743 19670 5752
rect 19628 5710 19656 5743
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19536 5494 19748 5522
rect 19444 5086 19564 5114
rect 19432 5024 19484 5030
rect 19536 5001 19564 5086
rect 19432 4966 19484 4972
rect 19522 4992 19578 5001
rect 19444 4622 19472 4966
rect 19522 4927 19578 4936
rect 19260 4554 19380 4570
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19248 4548 19380 4554
rect 19300 4542 19380 4548
rect 19248 4490 19300 4496
rect 18786 4448 18842 4457
rect 18786 4383 18842 4392
rect 19338 4448 19394 4457
rect 19338 4383 19394 4392
rect 19352 4010 19380 4383
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 19444 3602 19472 4558
rect 19536 4457 19564 4927
rect 19616 4480 19668 4486
rect 19522 4448 19578 4457
rect 19616 4422 19668 4428
rect 19522 4383 19578 4392
rect 19522 4312 19578 4321
rect 19522 4247 19578 4256
rect 19536 4214 19564 4247
rect 19524 4208 19576 4214
rect 19524 4150 19576 4156
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19444 3482 19472 3538
rect 19352 3454 19472 3482
rect 19352 3058 19380 3454
rect 19536 3398 19564 3878
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19628 3126 19656 4422
rect 19616 3120 19668 3126
rect 19616 3062 19668 3068
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19720 2938 19748 5494
rect 19812 3466 19840 6326
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 19904 5778 19932 6054
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19996 5556 20024 6412
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 20272 5953 20300 6326
rect 20364 6254 20392 8434
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20444 7744 20496 7750
rect 20548 7721 20576 8366
rect 20444 7686 20496 7692
rect 20534 7712 20590 7721
rect 20456 6866 20484 7686
rect 20534 7647 20590 7656
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20548 6497 20576 6734
rect 20640 6730 20668 8774
rect 20732 7818 20760 9862
rect 20824 9722 20852 11172
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20824 8634 20852 8842
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20824 7002 20852 7278
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20810 6896 20866 6905
rect 20810 6831 20866 6840
rect 20628 6724 20680 6730
rect 20628 6666 20680 6672
rect 20534 6488 20590 6497
rect 20534 6423 20590 6432
rect 20824 6390 20852 6831
rect 20628 6384 20680 6390
rect 20442 6352 20498 6361
rect 20442 6287 20498 6296
rect 20626 6352 20628 6361
rect 20812 6384 20864 6390
rect 20680 6352 20682 6361
rect 20812 6326 20864 6332
rect 20626 6287 20682 6296
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20258 5944 20314 5953
rect 20258 5879 20314 5888
rect 20272 5624 20300 5879
rect 20272 5596 20392 5624
rect 19904 5528 20024 5556
rect 19904 5352 19932 5528
rect 19994 5468 20302 5477
rect 19994 5466 20000 5468
rect 20056 5466 20080 5468
rect 20136 5466 20160 5468
rect 20216 5466 20240 5468
rect 20296 5466 20302 5468
rect 20056 5414 20058 5466
rect 20238 5414 20240 5466
rect 19994 5412 20000 5414
rect 20056 5412 20080 5414
rect 20136 5412 20160 5414
rect 20216 5412 20240 5414
rect 20296 5412 20302 5414
rect 19994 5403 20302 5412
rect 19904 5324 20024 5352
rect 19996 4690 20024 5324
rect 20364 5250 20392 5596
rect 20272 5222 20392 5250
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19904 3738 19932 4626
rect 20272 4486 20300 5222
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 19994 4380 20302 4389
rect 19994 4378 20000 4380
rect 20056 4378 20080 4380
rect 20136 4378 20160 4380
rect 20216 4378 20240 4380
rect 20296 4378 20302 4380
rect 20056 4326 20058 4378
rect 20238 4326 20240 4378
rect 19994 4324 20000 4326
rect 20056 4324 20080 4326
rect 20136 4324 20160 4326
rect 20216 4324 20240 4326
rect 20296 4324 20302 4326
rect 19994 4315 20302 4324
rect 20364 4078 20392 5034
rect 20456 4282 20484 6287
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20548 4758 20576 6122
rect 20824 6089 20852 6190
rect 20810 6080 20866 6089
rect 20810 6015 20866 6024
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20640 5710 20668 5850
rect 20812 5840 20864 5846
rect 20812 5782 20864 5788
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20824 5370 20852 5782
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20536 4752 20588 4758
rect 20536 4694 20588 4700
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20640 4010 20668 4558
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19800 3460 19852 3466
rect 19800 3402 19852 3408
rect 19904 3194 19932 3674
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 19994 3292 20302 3301
rect 19994 3290 20000 3292
rect 20056 3290 20080 3292
rect 20136 3290 20160 3292
rect 20216 3290 20240 3292
rect 20296 3290 20302 3292
rect 20056 3238 20058 3290
rect 20238 3238 20240 3290
rect 19994 3236 20000 3238
rect 20056 3236 20080 3238
rect 20136 3236 20160 3238
rect 20216 3236 20240 3238
rect 20296 3236 20302 3238
rect 19994 3227 20302 3236
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19260 2910 19748 2938
rect 19260 2774 19288 2910
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19430 2816 19486 2825
rect 19168 2746 19288 2774
rect 18694 2544 18750 2553
rect 18694 2479 18750 2488
rect 18420 2372 18472 2378
rect 18420 2314 18472 2320
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17868 2304 17920 2310
rect 19168 2281 19196 2746
rect 17868 2246 17920 2252
rect 19154 2272 19210 2281
rect 19154 2207 19210 2216
rect 16764 1828 16816 1834
rect 16764 1770 16816 1776
rect 16212 1556 16264 1562
rect 16212 1498 16264 1504
rect 15476 944 15528 950
rect 14108 870 14228 898
rect 15476 886 15528 892
rect 15936 944 15988 950
rect 15936 886 15988 892
rect 17408 944 17460 950
rect 17408 886 17460 892
rect 14108 762 14136 870
rect 14200 800 14228 870
rect 15488 800 15516 886
rect 17420 800 17448 886
rect 19352 800 19380 2790
rect 20824 2774 20852 3470
rect 20916 3126 20944 15370
rect 21100 15162 21128 17546
rect 21088 15156 21140 15162
rect 21008 15116 21088 15144
rect 21008 12288 21036 15116
rect 21088 15098 21140 15104
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21100 14346 21128 14758
rect 21284 14362 21312 20295
rect 21652 19854 21680 24754
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22284 22500 22336 22506
rect 22284 22442 22336 22448
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21732 20392 21784 20398
rect 21732 20334 21784 20340
rect 21744 19961 21772 20334
rect 21822 20088 21878 20097
rect 21822 20023 21878 20032
rect 21730 19952 21786 19961
rect 21730 19887 21732 19896
rect 21784 19887 21786 19896
rect 21732 19858 21784 19864
rect 21640 19848 21692 19854
rect 21640 19790 21692 19796
rect 21836 19718 21864 20023
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21376 18290 21404 19246
rect 21744 18970 21772 19450
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21744 17542 21772 18566
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21362 15192 21418 15201
rect 21362 15127 21418 15136
rect 21376 14958 21404 15127
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 21180 14340 21232 14346
rect 21284 14334 21496 14362
rect 21180 14282 21232 14288
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 21100 13734 21128 13942
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21100 12442 21128 13466
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 21008 12260 21128 12288
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 21008 9586 21036 12106
rect 21100 12102 21128 12260
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21086 9344 21142 9353
rect 21086 9279 21142 9288
rect 20994 9072 21050 9081
rect 20994 9007 21050 9016
rect 21008 8673 21036 9007
rect 20994 8664 21050 8673
rect 20994 8599 21050 8608
rect 20994 8528 21050 8537
rect 21100 8498 21128 9279
rect 20994 8463 21050 8472
rect 21088 8492 21140 8498
rect 21008 8430 21036 8463
rect 21088 8434 21140 8440
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 21192 8072 21220 14282
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21284 12850 21312 13330
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21376 12730 21404 13874
rect 21284 12702 21404 12730
rect 21284 12442 21312 12702
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21468 12374 21496 14334
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21560 12170 21588 16934
rect 21652 13938 21680 17002
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21640 12368 21692 12374
rect 21640 12310 21692 12316
rect 21652 12238 21680 12310
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 10742 21404 11494
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21284 9586 21312 10542
rect 21364 9988 21416 9994
rect 21364 9930 21416 9936
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21376 8265 21404 9930
rect 21468 8537 21496 12038
rect 21744 11762 21772 17478
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21836 15434 21864 16186
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21836 13530 21864 13738
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21928 12850 21956 20402
rect 22112 20058 22140 20470
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22204 19961 22232 19994
rect 22190 19952 22246 19961
rect 22190 19887 22246 19896
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 22020 19514 22048 19790
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22098 19544 22154 19553
rect 22008 19508 22060 19514
rect 22098 19479 22154 19488
rect 22008 19450 22060 19456
rect 22112 19242 22140 19479
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 22204 17762 22232 19654
rect 22296 19378 22324 22442
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22388 19922 22416 20198
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22296 18834 22324 19314
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22112 17734 22232 17762
rect 22296 17746 22324 18770
rect 22284 17740 22336 17746
rect 22112 17678 22140 17734
rect 22284 17682 22336 17688
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22296 16794 22324 17682
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22112 14550 22140 14894
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 22008 13252 22060 13258
rect 22008 13194 22060 13200
rect 22020 13025 22048 13194
rect 22006 13016 22062 13025
rect 22006 12951 22062 12960
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 22006 12064 22062 12073
rect 21836 11830 21864 12038
rect 22006 11999 22062 12008
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21652 11354 21680 11698
rect 21822 11384 21878 11393
rect 21640 11348 21692 11354
rect 21822 11319 21824 11328
rect 21640 11290 21692 11296
rect 21876 11319 21878 11328
rect 21824 11290 21876 11296
rect 21652 11234 21680 11290
rect 21652 11206 21864 11234
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21454 8528 21510 8537
rect 21560 8498 21588 9862
rect 21454 8463 21510 8472
rect 21548 8492 21600 8498
rect 21468 8294 21496 8463
rect 21548 8434 21600 8440
rect 21456 8288 21508 8294
rect 21362 8256 21418 8265
rect 21456 8230 21508 8236
rect 21362 8191 21418 8200
rect 21192 8044 21404 8072
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 21008 5137 21036 7414
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21100 7002 21128 7142
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 21192 6882 21220 7142
rect 21100 6854 21220 6882
rect 21100 6798 21128 6854
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 21100 5545 21128 5646
rect 21180 5636 21232 5642
rect 21180 5578 21232 5584
rect 21086 5536 21142 5545
rect 21086 5471 21142 5480
rect 20994 5128 21050 5137
rect 20994 5063 21050 5072
rect 20996 4208 21048 4214
rect 20996 4150 21048 4156
rect 20904 3120 20956 3126
rect 20904 3062 20956 3068
rect 20902 2952 20958 2961
rect 21008 2938 21036 4150
rect 21086 3904 21142 3913
rect 21086 3839 21142 3848
rect 21100 3466 21128 3839
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 20958 2910 21036 2938
rect 20902 2887 20958 2896
rect 20916 2854 20944 2887
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 19430 2751 19486 2760
rect 19444 2446 19472 2751
rect 20732 2746 20852 2774
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19994 2204 20302 2213
rect 19994 2202 20000 2204
rect 20056 2202 20080 2204
rect 20136 2202 20160 2204
rect 20216 2202 20240 2204
rect 20296 2202 20302 2204
rect 20056 2150 20058 2202
rect 20238 2150 20240 2202
rect 19994 2148 20000 2150
rect 20056 2148 20080 2150
rect 20136 2148 20160 2150
rect 20216 2148 20240 2150
rect 20296 2148 20302 2150
rect 19994 2139 20302 2148
rect 20732 1630 20760 2746
rect 21192 2650 21220 5578
rect 21376 5302 21404 8044
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21560 7546 21588 7686
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21456 7336 21508 7342
rect 21454 7304 21456 7313
rect 21508 7304 21510 7313
rect 21454 7239 21510 7248
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21284 4826 21312 5170
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21284 4486 21312 4762
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 21364 4072 21416 4078
rect 21362 4040 21364 4049
rect 21416 4040 21418 4049
rect 21362 3975 21418 3984
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 20720 1624 20772 1630
rect 20720 1566 20772 1572
rect 21100 950 21128 2314
rect 21088 944 21140 950
rect 21088 886 21140 892
rect 21284 800 21312 3334
rect 21468 3097 21496 6598
rect 21652 5642 21680 10066
rect 21744 9761 21772 10950
rect 21730 9752 21786 9761
rect 21730 9687 21786 9696
rect 21836 5930 21864 11206
rect 22020 9738 22048 11999
rect 22112 11830 22140 14486
rect 22204 13938 22232 15030
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22204 13734 22232 13874
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22204 13326 22232 13670
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22204 12782 22232 13126
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22190 11928 22246 11937
rect 22190 11863 22246 11872
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 21928 9710 22048 9738
rect 21928 8974 21956 9710
rect 22020 9030 22140 9058
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21914 8800 21970 8809
rect 22020 8786 22048 9030
rect 21970 8758 22048 8786
rect 21914 8735 21970 8744
rect 22006 7032 22062 7041
rect 22006 6967 22062 6976
rect 21914 5944 21970 5953
rect 21836 5902 21914 5930
rect 21914 5879 21970 5888
rect 21640 5636 21692 5642
rect 21640 5578 21692 5584
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 21652 4146 21680 5238
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21454 3088 21510 3097
rect 21454 3023 21510 3032
rect 21928 2825 21956 5879
rect 22020 4826 22048 6967
rect 22112 6322 22140 9030
rect 22204 8634 22232 11863
rect 22296 10810 22324 16458
rect 22388 16046 22416 19858
rect 22664 19310 22692 22918
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 22836 19984 22888 19990
rect 22834 19952 22836 19961
rect 22888 19952 22890 19961
rect 22834 19887 22890 19896
rect 22848 19553 22876 19887
rect 22834 19544 22890 19553
rect 22834 19479 22890 19488
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22756 18426 22784 18702
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22558 15464 22614 15473
rect 22558 15399 22614 15408
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 22388 12850 22416 13262
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22388 11898 22416 12650
rect 22480 12434 22508 13670
rect 22572 13258 22600 15399
rect 22560 13252 22612 13258
rect 22560 13194 22612 13200
rect 22664 12434 22692 18226
rect 22756 16454 22784 18362
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22848 17202 22876 18226
rect 22928 17876 22980 17882
rect 22928 17818 22980 17824
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22756 13326 22784 15846
rect 22940 15162 22968 17818
rect 23032 16658 23060 18566
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 22836 13524 22888 13530
rect 22836 13466 22888 13472
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 22848 13326 22876 13466
rect 23032 13433 23060 13466
rect 23018 13424 23074 13433
rect 23018 13359 23074 13368
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22848 12918 22876 13262
rect 22836 12912 22888 12918
rect 22836 12854 22888 12860
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 22480 12406 22600 12434
rect 22664 12406 22876 12434
rect 22572 12322 22600 12406
rect 22572 12294 22784 12322
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22560 12164 22612 12170
rect 22560 12106 22612 12112
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22572 11778 22600 12106
rect 22388 11750 22600 11778
rect 22664 11762 22692 12174
rect 22652 11756 22704 11762
rect 22388 11626 22416 11750
rect 22652 11698 22704 11704
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22376 11620 22428 11626
rect 22376 11562 22428 11568
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22282 9888 22338 9897
rect 22282 9823 22338 9832
rect 22296 9625 22324 9823
rect 22282 9616 22338 9625
rect 22282 9551 22338 9560
rect 22388 9178 22416 11562
rect 22480 11393 22508 11630
rect 22560 11552 22612 11558
rect 22756 11506 22784 12294
rect 22560 11494 22612 11500
rect 22466 11384 22522 11393
rect 22466 11319 22522 11328
rect 22572 9654 22600 11494
rect 22664 11478 22784 11506
rect 22664 11354 22692 11478
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22650 10432 22706 10441
rect 22650 10367 22706 10376
rect 22664 10062 22692 10367
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22204 8401 22232 8570
rect 22388 8480 22416 9114
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22480 8634 22508 8774
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22388 8452 22508 8480
rect 22190 8392 22246 8401
rect 22190 8327 22246 8336
rect 22374 8392 22430 8401
rect 22374 8327 22430 8336
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 22112 5953 22140 6122
rect 22204 6118 22232 7822
rect 22296 7721 22324 8026
rect 22282 7712 22338 7721
rect 22282 7647 22338 7656
rect 22296 6254 22324 7647
rect 22388 7410 22416 8327
rect 22480 7478 22508 8452
rect 22664 8294 22692 9658
rect 22742 9616 22798 9625
rect 22742 9551 22798 9560
rect 22756 9518 22784 9551
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22664 8266 22784 8294
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22468 7472 22520 7478
rect 22468 7414 22520 7420
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22374 6624 22430 6633
rect 22374 6559 22430 6568
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22098 5944 22154 5953
rect 22098 5879 22154 5888
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 22204 4758 22232 6054
rect 22296 5166 22324 6190
rect 22388 5642 22416 6559
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22466 6352 22522 6361
rect 22466 6287 22522 6296
rect 22480 6089 22508 6287
rect 22466 6080 22522 6089
rect 22466 6015 22522 6024
rect 22376 5636 22428 5642
rect 22376 5578 22428 5584
rect 22572 5574 22600 6394
rect 22560 5568 22612 5574
rect 22560 5510 22612 5516
rect 22374 5400 22430 5409
rect 22374 5335 22430 5344
rect 22388 5302 22416 5335
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 22466 5264 22522 5273
rect 22466 5199 22468 5208
rect 22520 5199 22522 5208
rect 22468 5170 22520 5176
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22192 4752 22244 4758
rect 22192 4694 22244 4700
rect 22296 4282 22324 5102
rect 22664 4690 22692 7686
rect 22756 7410 22784 8266
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 22756 7041 22784 7346
rect 22742 7032 22798 7041
rect 22742 6967 22798 6976
rect 22848 6458 22876 12406
rect 22940 11830 22968 12786
rect 23032 12170 23060 13359
rect 23124 12918 23152 20198
rect 23308 18306 23336 20334
rect 23386 18728 23442 18737
rect 23386 18663 23442 18672
rect 23400 18630 23428 18663
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23308 18290 23428 18306
rect 23308 18284 23440 18290
rect 23308 18278 23388 18284
rect 23388 18226 23440 18232
rect 23204 18216 23256 18222
rect 23256 18164 23336 18170
rect 23204 18158 23336 18164
rect 23216 18142 23336 18158
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 23216 16250 23244 16390
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23308 16130 23336 18142
rect 23400 17270 23428 18226
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 23216 16102 23336 16130
rect 23112 12912 23164 12918
rect 23112 12854 23164 12860
rect 23112 12436 23164 12442
rect 23112 12378 23164 12384
rect 23020 12164 23072 12170
rect 23020 12106 23072 12112
rect 22928 11824 22980 11830
rect 22928 11766 22980 11772
rect 23018 11248 23074 11257
rect 23018 11183 23074 11192
rect 22926 11112 22982 11121
rect 23032 11082 23060 11183
rect 22926 11047 22982 11056
rect 23020 11076 23072 11082
rect 22940 6730 22968 11047
rect 23020 11018 23072 11024
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22744 6316 22796 6322
rect 22744 6258 22796 6264
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22652 4072 22704 4078
rect 22652 4014 22704 4020
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22204 3126 22232 3878
rect 22572 3738 22600 4014
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 22664 3602 22692 4014
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22756 2990 22784 6258
rect 22848 4622 22876 6394
rect 23032 6186 23060 8366
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 23032 5914 23060 6122
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 23018 5400 23074 5409
rect 23018 5335 23074 5344
rect 23032 5302 23060 5335
rect 23020 5296 23072 5302
rect 23020 5238 23072 5244
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22940 4758 22968 5170
rect 22928 4752 22980 4758
rect 22928 4694 22980 4700
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 22940 3602 22968 4218
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 21914 2816 21970 2825
rect 21914 2751 21970 2760
rect 22020 2514 22048 2926
rect 23124 2774 23152 12378
rect 23216 12238 23244 16102
rect 23386 15872 23442 15881
rect 23386 15807 23442 15816
rect 23296 15088 23348 15094
rect 23400 15065 23428 15807
rect 23296 15030 23348 15036
rect 23386 15056 23442 15065
rect 23308 13682 23336 15030
rect 23386 14991 23442 15000
rect 23492 14006 23520 21422
rect 23584 21078 23612 26250
rect 23768 24750 23796 26794
rect 24755 26684 25063 26693
rect 24755 26682 24761 26684
rect 24817 26682 24841 26684
rect 24897 26682 24921 26684
rect 24977 26682 25001 26684
rect 25057 26682 25063 26684
rect 24817 26630 24819 26682
rect 24999 26630 25001 26682
rect 24755 26628 24761 26630
rect 24817 26628 24841 26630
rect 24897 26628 24921 26630
rect 24977 26628 25001 26630
rect 25057 26628 25063 26630
rect 24755 26619 25063 26628
rect 25148 26382 25176 28354
rect 26884 26784 26936 26790
rect 26884 26726 26936 26732
rect 26896 26586 26924 26726
rect 27356 26586 27384 28478
rect 28998 28354 29054 29154
rect 30286 28506 30342 29154
rect 32218 28506 32274 29154
rect 34150 28506 34206 29154
rect 36082 28506 36138 29154
rect 37370 28506 37426 29154
rect 39302 28506 39358 29154
rect 30286 28478 30604 28506
rect 30286 28354 30342 28478
rect 26884 26580 26936 26586
rect 26884 26522 26936 26528
rect 27344 26580 27396 26586
rect 27344 26522 27396 26528
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 25136 26376 25188 26382
rect 25136 26318 25188 26324
rect 24755 25596 25063 25605
rect 24755 25594 24761 25596
rect 24817 25594 24841 25596
rect 24897 25594 24921 25596
rect 24977 25594 25001 25596
rect 25057 25594 25063 25596
rect 24817 25542 24819 25594
rect 24999 25542 25001 25594
rect 24755 25540 24761 25542
rect 24817 25540 24841 25542
rect 24897 25540 24921 25542
rect 24977 25540 25001 25542
rect 25057 25540 25063 25542
rect 24755 25531 25063 25540
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 24950 24712 25006 24721
rect 23768 22094 23796 24686
rect 23860 24138 23888 24686
rect 24950 24647 24952 24656
rect 25004 24647 25006 24656
rect 24952 24618 25004 24624
rect 24755 24508 25063 24517
rect 24755 24506 24761 24508
rect 24817 24506 24841 24508
rect 24897 24506 24921 24508
rect 24977 24506 25001 24508
rect 25057 24506 25063 24508
rect 24817 24454 24819 24506
rect 24999 24454 25001 24506
rect 24755 24452 24761 24454
rect 24817 24452 24841 24454
rect 24897 24452 24921 24454
rect 24977 24452 25001 24454
rect 25057 24452 25063 24454
rect 24755 24443 25063 24452
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 25148 23798 25176 25230
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 24492 23656 24544 23662
rect 24492 23598 24544 23604
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 23768 22066 23888 22094
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23572 21072 23624 21078
rect 23572 21014 23624 21020
rect 23584 20806 23612 21014
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23676 20466 23704 21082
rect 23860 20466 23888 22066
rect 23664 20460 23716 20466
rect 23848 20460 23900 20466
rect 23716 20420 23796 20448
rect 23664 20402 23716 20408
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23570 20088 23626 20097
rect 23570 20023 23626 20032
rect 23584 16658 23612 20023
rect 23676 17678 23704 20198
rect 23768 18222 23796 20420
rect 23848 20402 23900 20408
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 23860 18034 23888 20402
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 23768 18006 23888 18034
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23662 17096 23718 17105
rect 23662 17031 23718 17040
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23584 16250 23612 16594
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23676 14346 23704 17031
rect 23768 16454 23796 18006
rect 23952 17338 23980 19382
rect 24136 19174 24164 22918
rect 24400 22772 24452 22778
rect 24400 22714 24452 22720
rect 24412 22642 24440 22714
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24124 19168 24176 19174
rect 24124 19110 24176 19116
rect 24032 18692 24084 18698
rect 24032 18634 24084 18640
rect 24044 18426 24072 18634
rect 24032 18420 24084 18426
rect 24032 18362 24084 18368
rect 24136 17338 24164 19110
rect 24504 18426 24532 23598
rect 24755 23420 25063 23429
rect 24755 23418 24761 23420
rect 24817 23418 24841 23420
rect 24897 23418 24921 23420
rect 24977 23418 25001 23420
rect 25057 23418 25063 23420
rect 24817 23366 24819 23418
rect 24999 23366 25001 23418
rect 24755 23364 24761 23366
rect 24817 23364 24841 23366
rect 24897 23364 24921 23366
rect 24977 23364 25001 23366
rect 25057 23364 25063 23366
rect 24755 23355 25063 23364
rect 24755 22332 25063 22341
rect 24755 22330 24761 22332
rect 24817 22330 24841 22332
rect 24897 22330 24921 22332
rect 24977 22330 25001 22332
rect 25057 22330 25063 22332
rect 24817 22278 24819 22330
rect 24999 22278 25001 22330
rect 24755 22276 24761 22278
rect 24817 22276 24841 22278
rect 24897 22276 24921 22278
rect 24977 22276 25001 22278
rect 25057 22276 25063 22278
rect 24755 22267 25063 22276
rect 25044 21956 25096 21962
rect 25044 21898 25096 21904
rect 25056 21486 25084 21898
rect 25148 21622 25176 23734
rect 25516 23118 25544 24754
rect 26976 24200 27028 24206
rect 26976 24142 27028 24148
rect 26424 23792 26476 23798
rect 26424 23734 26476 23740
rect 26240 23724 26292 23730
rect 26240 23666 26292 23672
rect 26252 23322 26280 23666
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 25320 23112 25372 23118
rect 25320 23054 25372 23060
rect 25504 23112 25556 23118
rect 25504 23054 25556 23060
rect 25228 22568 25280 22574
rect 25228 22510 25280 22516
rect 25240 22234 25268 22510
rect 25228 22228 25280 22234
rect 25228 22170 25280 22176
rect 25136 21616 25188 21622
rect 25136 21558 25188 21564
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 24755 21244 25063 21253
rect 24755 21242 24761 21244
rect 24817 21242 24841 21244
rect 24897 21242 24921 21244
rect 24977 21242 25001 21244
rect 25057 21242 25063 21244
rect 24817 21190 24819 21242
rect 24999 21190 25001 21242
rect 24755 21188 24761 21190
rect 24817 21188 24841 21190
rect 24897 21188 24921 21190
rect 24977 21188 25001 21190
rect 25057 21188 25063 21190
rect 24755 21179 25063 21188
rect 25148 21010 25176 21558
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 24596 19514 24624 20946
rect 25136 20324 25188 20330
rect 25136 20266 25188 20272
rect 24755 20156 25063 20165
rect 24755 20154 24761 20156
rect 24817 20154 24841 20156
rect 24897 20154 24921 20156
rect 24977 20154 25001 20156
rect 25057 20154 25063 20156
rect 24817 20102 24819 20154
rect 24999 20102 25001 20154
rect 24755 20100 24761 20102
rect 24817 20100 24841 20102
rect 24897 20100 24921 20102
rect 24977 20100 25001 20102
rect 25057 20100 25063 20102
rect 24755 20091 25063 20100
rect 24584 19508 24636 19514
rect 24584 19450 24636 19456
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24596 19378 24624 19450
rect 24780 19417 24808 19450
rect 24766 19408 24822 19417
rect 24584 19372 24636 19378
rect 24766 19343 24822 19352
rect 24584 19314 24636 19320
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 24596 17270 24624 19314
rect 24755 19068 25063 19077
rect 24755 19066 24761 19068
rect 24817 19066 24841 19068
rect 24897 19066 24921 19068
rect 24977 19066 25001 19068
rect 25057 19066 25063 19068
rect 24817 19014 24819 19066
rect 24999 19014 25001 19066
rect 24755 19012 24761 19014
rect 24817 19012 24841 19014
rect 24897 19012 24921 19014
rect 24977 19012 25001 19014
rect 25057 19012 25063 19014
rect 24755 19003 25063 19012
rect 25148 18834 25176 20266
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25148 18222 25176 18770
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 24755 17980 25063 17989
rect 24755 17978 24761 17980
rect 24817 17978 24841 17980
rect 24897 17978 24921 17980
rect 24977 17978 25001 17980
rect 25057 17978 25063 17980
rect 24817 17926 24819 17978
rect 24999 17926 25001 17978
rect 24755 17924 24761 17926
rect 24817 17924 24841 17926
rect 24897 17924 24921 17926
rect 24977 17924 25001 17926
rect 25057 17924 25063 17926
rect 24755 17915 25063 17924
rect 24950 17776 25006 17785
rect 24950 17711 25006 17720
rect 24964 17678 24992 17711
rect 24952 17672 25004 17678
rect 24674 17640 24730 17649
rect 24952 17614 25004 17620
rect 24674 17575 24730 17584
rect 24584 17264 24636 17270
rect 24584 17206 24636 17212
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 23860 16590 23888 17138
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23664 14340 23716 14346
rect 23664 14282 23716 14288
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 23308 13654 23428 13682
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23216 11665 23244 12174
rect 23202 11656 23258 11665
rect 23202 11591 23258 11600
rect 23204 10124 23256 10130
rect 23308 10112 23336 13194
rect 23256 10084 23336 10112
rect 23204 10066 23256 10072
rect 23216 5914 23244 10066
rect 23294 8120 23350 8129
rect 23294 8055 23350 8064
rect 23308 7886 23336 8055
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23400 7546 23428 13654
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23676 12442 23704 13126
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 23768 11150 23796 16390
rect 23860 15502 23888 16526
rect 24504 16522 24532 17138
rect 24492 16516 24544 16522
rect 24492 16458 24544 16464
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23952 15094 23980 15302
rect 23940 15088 23992 15094
rect 23940 15030 23992 15036
rect 24122 14920 24178 14929
rect 24122 14855 24178 14864
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23860 14006 23888 14214
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23860 12238 23888 13262
rect 23940 13184 23992 13190
rect 23940 13126 23992 13132
rect 23952 12617 23980 13126
rect 23938 12608 23994 12617
rect 23938 12543 23994 12552
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23952 11354 23980 11766
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 23756 11144 23808 11150
rect 23570 11112 23626 11121
rect 23756 11086 23808 11092
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23570 11047 23572 11056
rect 23624 11047 23626 11056
rect 23572 11018 23624 11024
rect 23480 8968 23532 8974
rect 23584 8956 23612 11018
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23676 9586 23704 10406
rect 23768 10062 23796 11086
rect 23860 10810 23888 11086
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 23756 10056 23808 10062
rect 23756 9998 23808 10004
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23676 9042 23704 9522
rect 23768 9450 23796 9862
rect 23756 9444 23808 9450
rect 23756 9386 23808 9392
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23532 8928 23612 8956
rect 23480 8910 23532 8916
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23296 7472 23348 7478
rect 23296 7414 23348 7420
rect 23308 6390 23336 7414
rect 23296 6384 23348 6390
rect 23296 6326 23348 6332
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23216 3602 23244 4558
rect 23204 3596 23256 3602
rect 23204 3538 23256 3544
rect 23400 3534 23428 4626
rect 23492 4554 23520 7890
rect 23676 6866 23704 8978
rect 23860 8634 23888 10746
rect 23952 9654 23980 10746
rect 23940 9648 23992 9654
rect 23940 9590 23992 9596
rect 24032 9648 24084 9654
rect 24032 9590 24084 9596
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 24044 8566 24072 9590
rect 24032 8560 24084 8566
rect 24032 8502 24084 8508
rect 23756 8016 23808 8022
rect 23940 8016 23992 8022
rect 23808 7976 23940 8004
rect 23756 7958 23808 7964
rect 23940 7958 23992 7964
rect 23940 7812 23992 7818
rect 23940 7754 23992 7760
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23754 7440 23810 7449
rect 23754 7375 23756 7384
rect 23808 7375 23810 7384
rect 23756 7346 23808 7352
rect 23860 7313 23888 7686
rect 23846 7304 23902 7313
rect 23846 7239 23902 7248
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23584 4622 23612 6190
rect 23848 5160 23900 5166
rect 23848 5102 23900 5108
rect 23860 5001 23888 5102
rect 23846 4992 23902 5001
rect 23846 4927 23902 4936
rect 23952 4758 23980 7754
rect 24136 7546 24164 14855
rect 24688 14521 24716 17575
rect 24755 16892 25063 16901
rect 24755 16890 24761 16892
rect 24817 16890 24841 16892
rect 24897 16890 24921 16892
rect 24977 16890 25001 16892
rect 25057 16890 25063 16892
rect 24817 16838 24819 16890
rect 24999 16838 25001 16890
rect 24755 16836 24761 16838
rect 24817 16836 24841 16838
rect 24897 16836 24921 16838
rect 24977 16836 25001 16838
rect 25057 16836 25063 16838
rect 24755 16827 25063 16836
rect 25148 16726 25176 18158
rect 25240 17746 25268 22170
rect 25332 18290 25360 23054
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25424 18834 25452 20538
rect 25516 20398 25544 23054
rect 26436 22953 26464 23734
rect 26516 23520 26568 23526
rect 26516 23462 26568 23468
rect 26422 22944 26478 22953
rect 26422 22879 26478 22888
rect 25596 20800 25648 20806
rect 25596 20742 25648 20748
rect 25504 20392 25556 20398
rect 25504 20334 25556 20340
rect 25516 18902 25544 20334
rect 25608 19718 25636 20742
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 25778 20088 25834 20097
rect 25778 20023 25834 20032
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25504 18896 25556 18902
rect 25504 18838 25556 18844
rect 25412 18828 25464 18834
rect 25412 18770 25464 18776
rect 25424 18698 25452 18770
rect 25412 18692 25464 18698
rect 25412 18634 25464 18640
rect 25424 18601 25452 18634
rect 25410 18592 25466 18601
rect 25410 18527 25466 18536
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25332 17785 25360 18226
rect 25318 17776 25374 17785
rect 25228 17740 25280 17746
rect 25318 17711 25374 17720
rect 25228 17682 25280 17688
rect 25136 16720 25188 16726
rect 25136 16662 25188 16668
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 24755 15804 25063 15813
rect 24755 15802 24761 15804
rect 24817 15802 24841 15804
rect 24897 15802 24921 15804
rect 24977 15802 25001 15804
rect 25057 15802 25063 15804
rect 24817 15750 24819 15802
rect 24999 15750 25001 15802
rect 24755 15748 24761 15750
rect 24817 15748 24841 15750
rect 24897 15748 24921 15750
rect 24977 15748 25001 15750
rect 25057 15748 25063 15750
rect 24755 15739 25063 15748
rect 24860 15632 24912 15638
rect 24858 15600 24860 15609
rect 24912 15600 24914 15609
rect 24858 15535 24914 15544
rect 25136 14952 25188 14958
rect 25134 14920 25136 14929
rect 25188 14920 25190 14929
rect 25134 14855 25190 14864
rect 24755 14716 25063 14725
rect 24755 14714 24761 14716
rect 24817 14714 24841 14716
rect 24897 14714 24921 14716
rect 24977 14714 25001 14716
rect 25057 14714 25063 14716
rect 24817 14662 24819 14714
rect 24999 14662 25001 14714
rect 24755 14660 24761 14662
rect 24817 14660 24841 14662
rect 24897 14660 24921 14662
rect 24977 14660 25001 14662
rect 25057 14660 25063 14662
rect 24755 14651 25063 14660
rect 24674 14512 24730 14521
rect 24674 14447 24730 14456
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24872 13938 24900 14418
rect 25240 14074 25268 16390
rect 25332 14482 25360 16594
rect 25504 15428 25556 15434
rect 25504 15370 25556 15376
rect 25320 14476 25372 14482
rect 25320 14418 25372 14424
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 24755 13628 25063 13637
rect 24755 13626 24761 13628
rect 24817 13626 24841 13628
rect 24897 13626 24921 13628
rect 24977 13626 25001 13628
rect 25057 13626 25063 13628
rect 24817 13574 24819 13626
rect 24999 13574 25001 13626
rect 24755 13572 24761 13574
rect 24817 13572 24841 13574
rect 24897 13572 24921 13574
rect 24977 13572 25001 13574
rect 25057 13572 25063 13574
rect 24755 13563 25063 13572
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24216 12708 24268 12714
rect 24216 12650 24268 12656
rect 24228 11014 24256 12650
rect 24504 12238 24532 12786
rect 24596 12434 24624 13262
rect 24755 12540 25063 12549
rect 24755 12538 24761 12540
rect 24817 12538 24841 12540
rect 24897 12538 24921 12540
rect 24977 12538 25001 12540
rect 25057 12538 25063 12540
rect 24817 12486 24819 12538
rect 24999 12486 25001 12538
rect 24755 12484 24761 12486
rect 24817 12484 24841 12486
rect 24897 12484 24921 12486
rect 24977 12484 25001 12486
rect 25057 12484 25063 12486
rect 24755 12475 25063 12484
rect 24596 12406 24716 12434
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24308 11076 24360 11082
rect 24308 11018 24360 11024
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24122 6624 24178 6633
rect 24122 6559 24178 6568
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24044 5030 24072 5102
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23480 4548 23532 4554
rect 23480 4490 23532 4496
rect 23848 4548 23900 4554
rect 23848 4490 23900 4496
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 23386 3360 23442 3369
rect 23386 3295 23442 3304
rect 23400 3058 23428 3295
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23124 2746 23244 2774
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 23216 2106 23244 2746
rect 23860 2582 23888 4490
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 24044 3534 24072 4082
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 24136 2990 24164 6559
rect 24228 6390 24256 10950
rect 24320 6905 24348 11018
rect 24504 10996 24532 12038
rect 24596 11150 24624 12174
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24504 10968 24624 10996
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24400 10532 24452 10538
rect 24400 10474 24452 10480
rect 24412 10130 24440 10474
rect 24504 10130 24532 10542
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24490 9616 24546 9625
rect 24490 9551 24546 9560
rect 24504 8906 24532 9551
rect 24492 8900 24544 8906
rect 24492 8842 24544 8848
rect 24400 8492 24452 8498
rect 24400 8434 24452 8440
rect 24306 6896 24362 6905
rect 24306 6831 24362 6840
rect 24216 6384 24268 6390
rect 24216 6326 24268 6332
rect 24412 4622 24440 8434
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 24412 3602 24440 4558
rect 24504 4282 24532 7346
rect 24596 7188 24624 10968
rect 24688 8809 24716 12406
rect 25148 12306 25176 13806
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 25148 11898 25176 12242
rect 25136 11892 25188 11898
rect 25136 11834 25188 11840
rect 24768 11824 24820 11830
rect 24766 11792 24768 11801
rect 24820 11792 24822 11801
rect 24766 11727 24822 11736
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 24755 11452 25063 11461
rect 24755 11450 24761 11452
rect 24817 11450 24841 11452
rect 24897 11450 24921 11452
rect 24977 11450 25001 11452
rect 25057 11450 25063 11452
rect 24817 11398 24819 11450
rect 24999 11398 25001 11450
rect 24755 11396 24761 11398
rect 24817 11396 24841 11398
rect 24897 11396 24921 11398
rect 24977 11396 25001 11398
rect 25057 11396 25063 11398
rect 24755 11387 25063 11396
rect 25148 11286 25176 11494
rect 25136 11280 25188 11286
rect 25136 11222 25188 11228
rect 24768 10736 24820 10742
rect 24766 10704 24768 10713
rect 24820 10704 24822 10713
rect 24766 10639 24822 10648
rect 25148 10606 25176 11222
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 25056 10452 25084 10542
rect 25056 10424 25176 10452
rect 24755 10364 25063 10373
rect 24755 10362 24761 10364
rect 24817 10362 24841 10364
rect 24897 10362 24921 10364
rect 24977 10362 25001 10364
rect 25057 10362 25063 10364
rect 24817 10310 24819 10362
rect 24999 10310 25001 10362
rect 24755 10308 24761 10310
rect 24817 10308 24841 10310
rect 24897 10308 24921 10310
rect 24977 10308 25001 10310
rect 25057 10308 25063 10310
rect 24755 10299 25063 10308
rect 25148 10305 25176 10424
rect 25134 10296 25190 10305
rect 25134 10231 25190 10240
rect 25044 10056 25096 10062
rect 24872 10016 25044 10044
rect 24872 10010 24900 10016
rect 24780 9994 24900 10010
rect 25044 9998 25096 10004
rect 24768 9988 24900 9994
rect 24820 9982 24900 9988
rect 24768 9930 24820 9936
rect 25044 9920 25096 9926
rect 25042 9888 25044 9897
rect 25096 9888 25098 9897
rect 25042 9823 25098 9832
rect 25134 9752 25190 9761
rect 25134 9687 25190 9696
rect 25148 9586 25176 9687
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 24755 9276 25063 9285
rect 24755 9274 24761 9276
rect 24817 9274 24841 9276
rect 24897 9274 24921 9276
rect 24977 9274 25001 9276
rect 25057 9274 25063 9276
rect 24817 9222 24819 9274
rect 24999 9222 25001 9274
rect 24755 9220 24761 9222
rect 24817 9220 24841 9222
rect 24897 9220 24921 9222
rect 24977 9220 25001 9222
rect 25057 9220 25063 9222
rect 24755 9211 25063 9220
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24674 8800 24730 8809
rect 24674 8735 24730 8744
rect 24872 8634 24900 8842
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24768 8560 24820 8566
rect 24688 8520 24768 8548
rect 24688 7818 24716 8520
rect 24768 8502 24820 8508
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 24755 8188 25063 8197
rect 24755 8186 24761 8188
rect 24817 8186 24841 8188
rect 24897 8186 24921 8188
rect 24977 8186 25001 8188
rect 25057 8186 25063 8188
rect 24817 8134 24819 8186
rect 24999 8134 25001 8186
rect 24755 8132 24761 8134
rect 24817 8132 24841 8134
rect 24897 8132 24921 8134
rect 24977 8132 25001 8134
rect 25057 8132 25063 8134
rect 24755 8123 25063 8132
rect 24766 7984 24822 7993
rect 24766 7919 24768 7928
rect 24820 7919 24822 7928
rect 24860 7948 24912 7954
rect 24768 7890 24820 7896
rect 24860 7890 24912 7896
rect 24676 7812 24728 7818
rect 24676 7754 24728 7760
rect 24872 7342 24900 7890
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 24964 7426 24992 7822
rect 25148 7818 25176 8230
rect 25240 7818 25268 14010
rect 25516 12986 25544 15370
rect 25608 13410 25636 19654
rect 25792 17882 25820 20023
rect 25870 19952 25926 19961
rect 25870 19887 25926 19896
rect 25884 18290 25912 19887
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 25976 17649 26004 20198
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26344 18834 26372 19994
rect 26422 19680 26478 19689
rect 26422 19615 26478 19624
rect 26436 18834 26464 19615
rect 26332 18828 26384 18834
rect 26332 18770 26384 18776
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 26528 18426 26556 23462
rect 26884 23044 26936 23050
rect 26884 22986 26936 22992
rect 26896 22574 26924 22986
rect 26884 22568 26936 22574
rect 26884 22510 26936 22516
rect 26988 22386 27016 24142
rect 26896 22358 27016 22386
rect 26700 22024 26752 22030
rect 26700 21966 26752 21972
rect 26608 18964 26660 18970
rect 26608 18906 26660 18912
rect 26516 18420 26568 18426
rect 26516 18362 26568 18368
rect 26620 18290 26648 18906
rect 26608 18284 26660 18290
rect 26608 18226 26660 18232
rect 26332 18216 26384 18222
rect 26054 18184 26110 18193
rect 26332 18158 26384 18164
rect 26054 18119 26056 18128
rect 26108 18119 26110 18128
rect 26056 18090 26108 18096
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 26160 17882 26188 18022
rect 26148 17876 26200 17882
rect 26148 17818 26200 17824
rect 25962 17640 26018 17649
rect 25962 17575 25964 17584
rect 26016 17575 26018 17584
rect 25964 17546 26016 17552
rect 26344 17338 26372 18158
rect 26332 17332 26384 17338
rect 26332 17274 26384 17280
rect 26712 17270 26740 21966
rect 26896 20602 26924 22358
rect 27448 22094 27476 26522
rect 27896 26444 27948 26450
rect 27896 26386 27948 26392
rect 27804 25356 27856 25362
rect 27804 25298 27856 25304
rect 27620 24608 27672 24614
rect 27620 24550 27672 24556
rect 27526 24168 27582 24177
rect 27526 24103 27528 24112
rect 27580 24103 27582 24112
rect 27528 24074 27580 24080
rect 27632 24070 27660 24550
rect 27712 24200 27764 24206
rect 27712 24142 27764 24148
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 27724 22098 27752 24142
rect 26988 22066 27476 22094
rect 27712 22092 27764 22098
rect 26884 20596 26936 20602
rect 26884 20538 26936 20544
rect 26988 20210 27016 22066
rect 27712 22034 27764 22040
rect 27618 21992 27674 22001
rect 27618 21927 27674 21936
rect 27632 21690 27660 21927
rect 27620 21684 27672 21690
rect 27620 21626 27672 21632
rect 27528 20392 27580 20398
rect 27528 20334 27580 20340
rect 26896 20182 27016 20210
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 26792 18828 26844 18834
rect 26792 18770 26844 18776
rect 26700 17264 26752 17270
rect 26606 17232 26662 17241
rect 26056 17196 26108 17202
rect 26700 17206 26752 17212
rect 26606 17167 26662 17176
rect 26056 17138 26108 17144
rect 26068 17105 26096 17138
rect 26054 17096 26110 17105
rect 26054 17031 26110 17040
rect 26620 16794 26648 17167
rect 26608 16788 26660 16794
rect 26608 16730 26660 16736
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25792 15434 25820 16594
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26422 16552 26478 16561
rect 26344 15502 26372 16526
rect 26422 16487 26478 16496
rect 26436 15706 26464 16487
rect 26700 16040 26752 16046
rect 26700 15982 26752 15988
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 25780 15428 25832 15434
rect 25780 15370 25832 15376
rect 25688 15360 25740 15366
rect 25686 15328 25688 15337
rect 25740 15328 25742 15337
rect 25686 15263 25742 15272
rect 26252 15094 26280 15438
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 25872 13728 25924 13734
rect 25872 13670 25924 13676
rect 25608 13382 25728 13410
rect 25596 13252 25648 13258
rect 25596 13194 25648 13200
rect 25504 12980 25556 12986
rect 25504 12922 25556 12928
rect 25504 12640 25556 12646
rect 25504 12582 25556 12588
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25424 11529 25452 12106
rect 25410 11520 25466 11529
rect 25410 11455 25466 11464
rect 25318 11384 25374 11393
rect 25318 11319 25374 11328
rect 25332 11121 25360 11319
rect 25318 11112 25374 11121
rect 25318 11047 25374 11056
rect 25424 10656 25452 11455
rect 25516 11098 25544 12582
rect 25608 12209 25636 13194
rect 25700 12646 25728 13382
rect 25884 13190 25912 13670
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 26160 12918 26188 13330
rect 26252 12986 26280 15030
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 25872 12844 25924 12850
rect 25872 12786 25924 12792
rect 25884 12646 25912 12786
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25594 12200 25650 12209
rect 25594 12135 25650 12144
rect 25608 11937 25636 12135
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25594 11928 25650 11937
rect 25594 11863 25650 11872
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 25608 11354 25636 11562
rect 25700 11558 25728 12038
rect 25780 11824 25832 11830
rect 25778 11792 25780 11801
rect 25832 11792 25834 11801
rect 25778 11727 25834 11736
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25688 11280 25740 11286
rect 25740 11240 25820 11268
rect 25688 11222 25740 11228
rect 25594 11112 25650 11121
rect 25516 11070 25594 11098
rect 25594 11047 25650 11056
rect 25608 11014 25636 11047
rect 25792 11014 25820 11240
rect 25596 11008 25648 11014
rect 25780 11008 25832 11014
rect 25596 10950 25648 10956
rect 25686 10976 25742 10985
rect 25780 10950 25832 10956
rect 25686 10911 25742 10920
rect 25596 10668 25648 10674
rect 25424 10628 25544 10656
rect 25410 10568 25466 10577
rect 25410 10503 25466 10512
rect 25318 10432 25374 10441
rect 25318 10367 25374 10376
rect 25332 9654 25360 10367
rect 25424 9897 25452 10503
rect 25516 10470 25544 10628
rect 25596 10610 25648 10616
rect 25608 10577 25636 10610
rect 25594 10568 25650 10577
rect 25594 10503 25650 10512
rect 25504 10464 25556 10470
rect 25596 10464 25648 10470
rect 25504 10406 25556 10412
rect 25594 10432 25596 10441
rect 25648 10432 25650 10441
rect 25594 10367 25650 10376
rect 25596 10192 25648 10198
rect 25596 10134 25648 10140
rect 25410 9888 25466 9897
rect 25410 9823 25466 9832
rect 25320 9648 25372 9654
rect 25320 9590 25372 9596
rect 25332 9382 25360 9590
rect 25608 9382 25636 10134
rect 25700 9994 25728 10911
rect 25884 10826 25912 12582
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 25976 11762 26004 12242
rect 26068 11898 26096 12378
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 26068 11336 26096 11834
rect 26160 11694 26188 12854
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 26252 11801 26280 12786
rect 26238 11792 26294 11801
rect 26238 11727 26294 11736
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 26240 11620 26292 11626
rect 26240 11562 26292 11568
rect 25792 10798 25912 10826
rect 25976 11308 26096 11336
rect 26146 11384 26202 11393
rect 26146 11319 26202 11328
rect 25976 10810 26004 11308
rect 26056 11212 26108 11218
rect 26056 11154 26108 11160
rect 25964 10804 26016 10810
rect 25688 9988 25740 9994
rect 25688 9930 25740 9936
rect 25688 9580 25740 9586
rect 25688 9522 25740 9528
rect 25320 9376 25372 9382
rect 25504 9376 25556 9382
rect 25320 9318 25372 9324
rect 25410 9344 25466 9353
rect 25504 9318 25556 9324
rect 25596 9376 25648 9382
rect 25596 9318 25648 9324
rect 25410 9279 25466 9288
rect 25318 9208 25374 9217
rect 25318 9143 25374 9152
rect 25136 7812 25188 7818
rect 25136 7754 25188 7760
rect 25228 7812 25280 7818
rect 25228 7754 25280 7760
rect 25332 7750 25360 9143
rect 25424 8242 25452 9279
rect 25516 8362 25544 9318
rect 25608 9178 25636 9318
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25594 8528 25650 8537
rect 25594 8463 25650 8472
rect 25608 8430 25636 8463
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 25700 8362 25728 9522
rect 25792 8498 25820 10798
rect 25964 10746 26016 10752
rect 25870 10432 25926 10441
rect 25870 10367 25926 10376
rect 25884 9926 25912 10367
rect 25872 9920 25924 9926
rect 25872 9862 25924 9868
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25504 8356 25556 8362
rect 25504 8298 25556 8304
rect 25688 8356 25740 8362
rect 25688 8298 25740 8304
rect 25424 8214 25728 8242
rect 25504 7812 25556 7818
rect 25504 7754 25556 7760
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25516 7478 25544 7754
rect 25596 7744 25648 7750
rect 25596 7686 25648 7692
rect 25228 7472 25280 7478
rect 25042 7440 25098 7449
rect 24964 7398 25042 7426
rect 25504 7472 25556 7478
rect 25228 7414 25280 7420
rect 25318 7440 25374 7449
rect 25042 7375 25098 7384
rect 24860 7336 24912 7342
rect 24860 7278 24912 7284
rect 25136 7336 25188 7342
rect 25240 7313 25268 7414
rect 25318 7375 25374 7384
rect 25502 7440 25504 7449
rect 25556 7440 25558 7449
rect 25502 7375 25558 7384
rect 25136 7278 25188 7284
rect 25226 7304 25282 7313
rect 24860 7200 24912 7206
rect 24596 7160 24860 7188
rect 24596 5914 24624 7160
rect 24860 7142 24912 7148
rect 24755 7100 25063 7109
rect 24755 7098 24761 7100
rect 24817 7098 24841 7100
rect 24897 7098 24921 7100
rect 24977 7098 25001 7100
rect 25057 7098 25063 7100
rect 24817 7046 24819 7098
rect 24999 7046 25001 7098
rect 24755 7044 24761 7046
rect 24817 7044 24841 7046
rect 24897 7044 24921 7046
rect 24977 7044 25001 7046
rect 25057 7044 25063 7046
rect 24755 7035 25063 7044
rect 25148 6866 25176 7278
rect 25226 7239 25282 7248
rect 25332 7177 25360 7375
rect 25318 7168 25374 7177
rect 25318 7103 25374 7112
rect 25226 7032 25282 7041
rect 25226 6967 25228 6976
rect 25280 6967 25282 6976
rect 25228 6938 25280 6944
rect 25332 6866 25452 6882
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25332 6860 25464 6866
rect 25332 6854 25412 6860
rect 25332 6769 25360 6854
rect 25412 6802 25464 6808
rect 25318 6760 25374 6769
rect 25318 6695 25374 6704
rect 25412 6724 25464 6730
rect 24768 6384 24820 6390
rect 24768 6326 24820 6332
rect 24780 6118 24808 6326
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24755 6012 25063 6021
rect 24755 6010 24761 6012
rect 24817 6010 24841 6012
rect 24897 6010 24921 6012
rect 24977 6010 25001 6012
rect 25057 6010 25063 6012
rect 24817 5958 24819 6010
rect 24999 5958 25001 6010
rect 24755 5956 24761 5958
rect 24817 5956 24841 5958
rect 24897 5956 24921 5958
rect 24977 5956 25001 5958
rect 25057 5956 25063 5958
rect 24755 5947 25063 5956
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 25148 5778 25176 6190
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 24766 5672 24822 5681
rect 24766 5607 24768 5616
rect 24820 5607 24822 5616
rect 24768 5578 24820 5584
rect 25148 5302 25176 5714
rect 25332 5710 25360 6695
rect 25412 6666 25464 6672
rect 25424 5914 25452 6666
rect 25516 6390 25544 7375
rect 25504 6384 25556 6390
rect 25504 6326 25556 6332
rect 25608 6066 25636 7686
rect 25700 7546 25728 8214
rect 25884 7886 25912 9862
rect 25976 9353 26004 10746
rect 25962 9344 26018 9353
rect 25962 9279 26018 9288
rect 25962 9072 26018 9081
rect 25962 9007 26018 9016
rect 25976 8634 26004 9007
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 25976 8362 26004 8570
rect 25964 8356 26016 8362
rect 25964 8298 26016 8304
rect 26068 7993 26096 11154
rect 26160 9994 26188 11319
rect 26252 11150 26280 11562
rect 26344 11354 26372 14758
rect 26516 13728 26568 13734
rect 26516 13670 26568 13676
rect 26528 13190 26556 13670
rect 26620 13394 26648 15506
rect 26712 15434 26740 15982
rect 26700 15428 26752 15434
rect 26700 15370 26752 15376
rect 26804 15026 26832 18770
rect 26896 18698 26924 20182
rect 27172 19310 27200 20198
rect 27540 19514 27568 20334
rect 27528 19508 27580 19514
rect 27528 19450 27580 19456
rect 27160 19304 27212 19310
rect 27160 19246 27212 19252
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 26884 18692 26936 18698
rect 26884 18634 26936 18640
rect 26896 17610 26924 18634
rect 26976 18080 27028 18086
rect 27080 18057 27108 18838
rect 27724 18714 27752 22034
rect 27816 21146 27844 25298
rect 27908 23186 27936 26386
rect 29012 26382 29040 28354
rect 29182 26480 29238 26489
rect 29182 26415 29184 26424
rect 29236 26415 29238 26424
rect 29184 26386 29236 26392
rect 30576 26382 30604 28478
rect 32218 28478 32536 28506
rect 32218 28354 32274 28478
rect 32508 26586 32536 28478
rect 34150 28478 34652 28506
rect 34150 28354 34206 28478
rect 34152 26784 34204 26790
rect 34152 26726 34204 26732
rect 32496 26580 32548 26586
rect 32496 26522 32548 26528
rect 33600 26580 33652 26586
rect 33600 26522 33652 26528
rect 28632 26376 28684 26382
rect 28368 26336 28632 26364
rect 28264 26308 28316 26314
rect 28264 26250 28316 26256
rect 28172 24948 28224 24954
rect 28172 24890 28224 24896
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28092 24206 28120 24754
rect 28184 24410 28212 24890
rect 28172 24404 28224 24410
rect 28172 24346 28224 24352
rect 28080 24200 28132 24206
rect 28080 24142 28132 24148
rect 27896 23180 27948 23186
rect 27896 23122 27948 23128
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27816 18970 27844 20878
rect 27908 19310 27936 23122
rect 28276 22710 28304 26250
rect 28264 22704 28316 22710
rect 28264 22646 28316 22652
rect 28000 21010 28212 21026
rect 28000 21004 28224 21010
rect 28000 20998 28172 21004
rect 27896 19304 27948 19310
rect 27896 19246 27948 19252
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 27632 18686 27752 18714
rect 27908 18698 27936 19246
rect 27896 18692 27948 18698
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27172 18290 27200 18566
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 26976 18022 27028 18028
rect 27066 18048 27122 18057
rect 26884 17604 26936 17610
rect 26884 17546 26936 17552
rect 26792 15020 26844 15026
rect 26792 14962 26844 14968
rect 26792 14612 26844 14618
rect 26792 14554 26844 14560
rect 26804 14362 26832 14554
rect 26712 14334 26832 14362
rect 26712 14278 26740 14334
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26804 13841 26832 14214
rect 26790 13832 26846 13841
rect 26790 13767 26846 13776
rect 26608 13388 26660 13394
rect 26608 13330 26660 13336
rect 26620 13274 26648 13330
rect 26620 13246 26740 13274
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26528 12986 26556 13126
rect 26516 12980 26568 12986
rect 26516 12922 26568 12928
rect 26608 12776 26660 12782
rect 26608 12718 26660 12724
rect 26620 12322 26648 12718
rect 26712 12442 26740 13246
rect 26792 13252 26844 13258
rect 26792 13194 26844 13200
rect 26804 12889 26832 13194
rect 26790 12880 26846 12889
rect 26790 12815 26846 12824
rect 26896 12764 26924 17546
rect 26804 12736 26924 12764
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 26620 12294 26740 12322
rect 26424 11824 26476 11830
rect 26424 11766 26476 11772
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 26436 11218 26464 11766
rect 26608 11348 26660 11354
rect 26528 11308 26608 11336
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26424 11076 26476 11082
rect 26424 11018 26476 11024
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26252 10470 26280 10610
rect 26240 10464 26292 10470
rect 26240 10406 26292 10412
rect 26148 9988 26200 9994
rect 26148 9930 26200 9936
rect 26240 9920 26292 9926
rect 26240 9862 26292 9868
rect 26148 9444 26200 9450
rect 26148 9386 26200 9392
rect 26054 7984 26110 7993
rect 26054 7919 26056 7928
rect 26108 7919 26110 7928
rect 26056 7890 26108 7896
rect 25872 7880 25924 7886
rect 25872 7822 25924 7828
rect 25964 7812 26016 7818
rect 25964 7754 26016 7760
rect 26056 7812 26108 7818
rect 26056 7754 26108 7760
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 25780 7268 25832 7274
rect 25780 7210 25832 7216
rect 25792 6322 25820 7210
rect 25780 6316 25832 6322
rect 25780 6258 25832 6264
rect 25516 6038 25636 6066
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25320 5704 25372 5710
rect 25320 5646 25372 5652
rect 25136 5296 25188 5302
rect 25516 5273 25544 6038
rect 25594 5944 25650 5953
rect 25594 5879 25650 5888
rect 25608 5778 25636 5879
rect 25596 5772 25648 5778
rect 25596 5714 25648 5720
rect 25884 5574 25912 7482
rect 25976 7410 26004 7754
rect 26068 7721 26096 7754
rect 26054 7712 26110 7721
rect 26054 7647 26110 7656
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25976 7206 26004 7346
rect 25964 7200 26016 7206
rect 25964 7142 26016 7148
rect 26160 7002 26188 9386
rect 26252 9178 26280 9862
rect 26240 9172 26292 9178
rect 26240 9114 26292 9120
rect 26252 8634 26280 9114
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 26344 7834 26372 10610
rect 26436 9178 26464 11018
rect 26528 10198 26556 11308
rect 26608 11290 26660 11296
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26516 10192 26568 10198
rect 26516 10134 26568 10140
rect 26620 10044 26648 11154
rect 26712 10606 26740 12294
rect 26804 11082 26832 12736
rect 26988 12617 27016 18022
rect 27066 17983 27122 17992
rect 27540 17921 27568 18566
rect 27526 17912 27582 17921
rect 27632 17882 27660 18686
rect 27896 18634 27948 18640
rect 28000 18578 28028 20998
rect 28172 20946 28224 20952
rect 28276 20806 28304 22646
rect 28172 20800 28224 20806
rect 28172 20742 28224 20748
rect 28264 20800 28316 20806
rect 28264 20742 28316 20748
rect 28184 19514 28212 20742
rect 28172 19508 28224 19514
rect 28172 19450 28224 19456
rect 28368 19417 28396 26336
rect 28632 26318 28684 26324
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 31116 26308 31168 26314
rect 31116 26250 31168 26256
rect 32404 26308 32456 26314
rect 32404 26250 32456 26256
rect 29516 26140 29824 26149
rect 29516 26138 29522 26140
rect 29578 26138 29602 26140
rect 29658 26138 29682 26140
rect 29738 26138 29762 26140
rect 29818 26138 29824 26140
rect 29578 26086 29580 26138
rect 29760 26086 29762 26138
rect 29516 26084 29522 26086
rect 29578 26084 29602 26086
rect 29658 26084 29682 26086
rect 29738 26084 29762 26086
rect 29818 26084 29824 26086
rect 29516 26075 29824 26084
rect 30196 25968 30248 25974
rect 30196 25910 30248 25916
rect 30208 25362 30236 25910
rect 30288 25900 30340 25906
rect 30288 25842 30340 25848
rect 30196 25356 30248 25362
rect 30196 25298 30248 25304
rect 28448 25152 28500 25158
rect 28448 25094 28500 25100
rect 28816 25152 28868 25158
rect 28816 25094 28868 25100
rect 28460 20874 28488 25094
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28552 22030 28580 24142
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28724 22024 28776 22030
rect 28724 21966 28776 21972
rect 28632 21888 28684 21894
rect 28632 21830 28684 21836
rect 28644 21622 28672 21830
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28552 20602 28580 21422
rect 28736 21146 28764 21966
rect 28724 21140 28776 21146
rect 28724 21082 28776 21088
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 28354 19408 28410 19417
rect 28354 19343 28410 19352
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 27724 18550 28028 18578
rect 27724 18222 27752 18550
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27526 17847 27582 17856
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27160 17808 27212 17814
rect 27160 17750 27212 17756
rect 27172 16998 27200 17750
rect 27344 17740 27396 17746
rect 27344 17682 27396 17688
rect 27252 17672 27304 17678
rect 27252 17614 27304 17620
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 27066 16688 27122 16697
rect 27066 16623 27122 16632
rect 26974 12608 27030 12617
rect 26974 12543 27030 12552
rect 26976 12096 27028 12102
rect 26976 12038 27028 12044
rect 26884 11620 26936 11626
rect 26884 11562 26936 11568
rect 26896 11150 26924 11562
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26792 11076 26844 11082
rect 26792 11018 26844 11024
rect 26884 11008 26936 11014
rect 26884 10950 26936 10956
rect 26700 10600 26752 10606
rect 26700 10542 26752 10548
rect 26790 10432 26846 10441
rect 26790 10367 26846 10376
rect 26804 10130 26832 10367
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26528 10016 26648 10044
rect 26528 9722 26556 10016
rect 26516 9716 26568 9722
rect 26516 9658 26568 9664
rect 26792 9648 26844 9654
rect 26792 9590 26844 9596
rect 26700 9580 26752 9586
rect 26700 9522 26752 9528
rect 26516 9444 26568 9450
rect 26516 9386 26568 9392
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26436 8838 26464 8978
rect 26424 8832 26476 8838
rect 26424 8774 26476 8780
rect 26528 8430 26556 9386
rect 26608 9172 26660 9178
rect 26608 9114 26660 9120
rect 26620 9042 26648 9114
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 26424 7948 26476 7954
rect 26424 7890 26476 7896
rect 26252 7806 26372 7834
rect 26148 6996 26200 7002
rect 26148 6938 26200 6944
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26056 5840 26108 5846
rect 26056 5782 26108 5788
rect 25964 5772 26016 5778
rect 25964 5714 26016 5720
rect 25872 5568 25924 5574
rect 25872 5510 25924 5516
rect 25136 5238 25188 5244
rect 25502 5264 25558 5273
rect 24676 5228 24728 5234
rect 25502 5199 25558 5208
rect 24676 5170 24728 5176
rect 24492 4276 24544 4282
rect 24492 4218 24544 4224
rect 24688 4010 24716 5170
rect 25778 4992 25834 5001
rect 24755 4924 25063 4933
rect 25778 4927 25834 4936
rect 24755 4922 24761 4924
rect 24817 4922 24841 4924
rect 24897 4922 24921 4924
rect 24977 4922 25001 4924
rect 25057 4922 25063 4924
rect 24817 4870 24819 4922
rect 24999 4870 25001 4922
rect 24755 4868 24761 4870
rect 24817 4868 24841 4870
rect 24897 4868 24921 4870
rect 24977 4868 25001 4870
rect 25057 4868 25063 4870
rect 24755 4859 25063 4868
rect 25792 4826 25820 4927
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 24768 4548 24820 4554
rect 24768 4490 24820 4496
rect 25780 4548 25832 4554
rect 25780 4490 25832 4496
rect 24780 4128 24808 4490
rect 24860 4140 24912 4146
rect 24780 4100 24860 4128
rect 24860 4082 24912 4088
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 24676 4004 24728 4010
rect 24676 3946 24728 3952
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24400 3596 24452 3602
rect 24320 3556 24400 3584
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 24320 2854 24348 3556
rect 24400 3538 24452 3544
rect 24308 2848 24360 2854
rect 24308 2790 24360 2796
rect 24504 2650 24532 3878
rect 24688 3602 24716 3946
rect 25148 3913 25176 4014
rect 25688 3936 25740 3942
rect 25134 3904 25190 3913
rect 25688 3878 25740 3884
rect 24755 3836 25063 3845
rect 25134 3839 25190 3848
rect 24755 3834 24761 3836
rect 24817 3834 24841 3836
rect 24897 3834 24921 3836
rect 24977 3834 25001 3836
rect 25057 3834 25063 3836
rect 24817 3782 24819 3834
rect 24999 3782 25001 3834
rect 24755 3780 24761 3782
rect 24817 3780 24841 3782
rect 24897 3780 24921 3782
rect 24977 3780 25001 3782
rect 25057 3780 25063 3782
rect 24755 3771 25063 3780
rect 25700 3738 25728 3878
rect 25688 3732 25740 3738
rect 25688 3674 25740 3680
rect 24676 3596 24728 3602
rect 24596 3556 24676 3584
rect 24596 3126 24624 3556
rect 24676 3538 24728 3544
rect 24584 3120 24636 3126
rect 24584 3062 24636 3068
rect 24492 2644 24544 2650
rect 24492 2586 24544 2592
rect 23848 2576 23900 2582
rect 23848 2518 23900 2524
rect 24596 2514 24624 3062
rect 25792 3058 25820 4490
rect 25976 3913 26004 5714
rect 26068 4826 26096 5782
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 26054 4040 26110 4049
rect 26160 4026 26188 6258
rect 26252 6118 26280 7806
rect 26332 7744 26384 7750
rect 26436 7721 26464 7890
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26332 7686 26384 7692
rect 26422 7712 26478 7721
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 26344 5914 26372 7686
rect 26422 7647 26478 7656
rect 26620 6934 26648 7822
rect 26608 6928 26660 6934
rect 26712 6905 26740 9522
rect 26804 9382 26832 9590
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26792 8968 26844 8974
rect 26792 8910 26844 8916
rect 26804 8430 26832 8910
rect 26792 8424 26844 8430
rect 26792 8366 26844 8372
rect 26804 7886 26832 8366
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26804 7342 26832 7822
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26608 6870 26660 6876
rect 26698 6896 26754 6905
rect 26516 6180 26568 6186
rect 26516 6122 26568 6128
rect 26422 5944 26478 5953
rect 26332 5908 26384 5914
rect 26422 5879 26478 5888
rect 26332 5850 26384 5856
rect 26436 5846 26464 5879
rect 26424 5840 26476 5846
rect 26424 5782 26476 5788
rect 26330 4720 26386 4729
rect 26330 4655 26386 4664
rect 26344 4622 26372 4655
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26240 4548 26292 4554
rect 26240 4490 26292 4496
rect 26252 4282 26280 4490
rect 26330 4448 26386 4457
rect 26330 4383 26386 4392
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 26240 4072 26292 4078
rect 26160 4020 26240 4026
rect 26160 4014 26292 4020
rect 26160 3998 26280 4014
rect 26054 3975 26110 3984
rect 25962 3904 26018 3913
rect 25962 3839 26018 3848
rect 26068 3126 26096 3975
rect 26148 3528 26200 3534
rect 26146 3496 26148 3505
rect 26200 3496 26202 3505
rect 26146 3431 26202 3440
rect 26056 3120 26108 3126
rect 26056 3062 26108 3068
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 24860 2984 24912 2990
rect 24688 2944 24860 2972
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24584 2372 24636 2378
rect 24584 2314 24636 2320
rect 23204 2100 23256 2106
rect 23204 2042 23256 2048
rect 24596 1834 24624 2314
rect 24584 1828 24636 1834
rect 24584 1770 24636 1776
rect 24688 1578 24716 2944
rect 24860 2926 24912 2932
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 24755 2748 25063 2757
rect 24755 2746 24761 2748
rect 24817 2746 24841 2748
rect 24897 2746 24921 2748
rect 24977 2746 25001 2748
rect 25057 2746 25063 2748
rect 24817 2694 24819 2746
rect 24999 2694 25001 2746
rect 24755 2692 24761 2694
rect 24817 2692 24841 2694
rect 24897 2692 24921 2694
rect 24977 2692 25001 2694
rect 25057 2692 25063 2694
rect 24755 2683 25063 2692
rect 25134 2680 25190 2689
rect 25134 2615 25190 2624
rect 25148 2378 25176 2615
rect 25318 2544 25374 2553
rect 25318 2479 25374 2488
rect 25332 2378 25360 2479
rect 25136 2372 25188 2378
rect 25136 2314 25188 2320
rect 25320 2372 25372 2378
rect 25320 2314 25372 2320
rect 25516 1698 25544 2858
rect 26344 2650 26372 4383
rect 26528 2774 26556 6122
rect 26620 4214 26648 6870
rect 26698 6831 26754 6840
rect 26712 5642 26740 6831
rect 26896 5778 26924 10950
rect 26988 7546 27016 12038
rect 27080 10674 27108 16623
rect 27172 11286 27200 16934
rect 27264 13954 27292 17614
rect 27356 16590 27384 17682
rect 27436 17536 27488 17542
rect 27436 17478 27488 17484
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 27448 17270 27476 17478
rect 27436 17264 27488 17270
rect 27436 17206 27488 17212
rect 27344 16584 27396 16590
rect 27344 16526 27396 16532
rect 27356 16114 27384 16526
rect 27540 16250 27568 17478
rect 27632 16998 27660 17818
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 27620 16516 27672 16522
rect 27620 16458 27672 16464
rect 27528 16244 27580 16250
rect 27528 16186 27580 16192
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27632 15706 27660 16458
rect 27620 15700 27672 15706
rect 27620 15642 27672 15648
rect 27620 14476 27672 14482
rect 27620 14418 27672 14424
rect 27264 13926 27384 13954
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27264 12170 27292 13806
rect 27356 12238 27384 13926
rect 27436 13932 27488 13938
rect 27436 13874 27488 13880
rect 27448 13462 27476 13874
rect 27436 13456 27488 13462
rect 27436 13398 27488 13404
rect 27448 12646 27476 13398
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 27252 12164 27304 12170
rect 27252 12106 27304 12112
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27160 11280 27212 11286
rect 27160 11222 27212 11228
rect 27160 11008 27212 11014
rect 27160 10950 27212 10956
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 27172 10538 27200 10950
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27160 10532 27212 10538
rect 27160 10474 27212 10480
rect 27160 10192 27212 10198
rect 27080 10152 27160 10180
rect 27080 7585 27108 10152
rect 27160 10134 27212 10140
rect 27160 9988 27212 9994
rect 27160 9930 27212 9936
rect 27172 9761 27200 9930
rect 27158 9752 27214 9761
rect 27158 9687 27214 9696
rect 27160 9444 27212 9450
rect 27160 9386 27212 9392
rect 27066 7576 27122 7585
rect 26976 7540 27028 7546
rect 27066 7511 27122 7520
rect 26976 7482 27028 7488
rect 27172 7002 27200 9386
rect 26976 6996 27028 7002
rect 26976 6938 27028 6944
rect 27160 6996 27212 7002
rect 27160 6938 27212 6944
rect 26884 5772 26936 5778
rect 26884 5714 26936 5720
rect 26792 5704 26844 5710
rect 26792 5646 26844 5652
rect 26700 5636 26752 5642
rect 26700 5578 26752 5584
rect 26804 5137 26832 5646
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 26790 5128 26846 5137
rect 26790 5063 26846 5072
rect 26608 4208 26660 4214
rect 26608 4150 26660 4156
rect 26608 3460 26660 3466
rect 26608 3402 26660 3408
rect 26620 3233 26648 3402
rect 26606 3224 26662 3233
rect 26606 3159 26662 3168
rect 26436 2746 26556 2774
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 25504 1692 25556 1698
rect 25504 1634 25556 1640
rect 24504 1550 24716 1578
rect 22560 944 22612 950
rect 22560 886 22612 892
rect 22572 800 22600 886
rect 24504 800 24532 1550
rect 26436 800 26464 2746
rect 26896 2650 26924 5238
rect 26988 5166 27016 6938
rect 27068 5772 27120 5778
rect 27068 5714 27120 5720
rect 26976 5160 27028 5166
rect 26976 5102 27028 5108
rect 27080 3194 27108 5714
rect 27264 4690 27292 10542
rect 27356 9926 27384 12038
rect 27448 10674 27476 12378
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27540 11830 27568 12038
rect 27528 11824 27580 11830
rect 27528 11766 27580 11772
rect 27528 11280 27580 11286
rect 27526 11248 27528 11257
rect 27580 11248 27582 11257
rect 27526 11183 27582 11192
rect 27526 10840 27582 10849
rect 27526 10775 27582 10784
rect 27436 10668 27488 10674
rect 27436 10610 27488 10616
rect 27434 10432 27490 10441
rect 27434 10367 27490 10376
rect 27448 10169 27476 10367
rect 27434 10160 27490 10169
rect 27434 10095 27490 10104
rect 27448 9994 27476 10095
rect 27540 9994 27568 10775
rect 27632 10198 27660 14418
rect 27724 13394 27752 18158
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 28000 14550 28028 16934
rect 28172 15632 28224 15638
rect 28092 15592 28172 15620
rect 27804 14544 27856 14550
rect 27804 14486 27856 14492
rect 27988 14544 28040 14550
rect 27988 14486 28040 14492
rect 27712 13388 27764 13394
rect 27712 13330 27764 13336
rect 27712 11076 27764 11082
rect 27712 11018 27764 11024
rect 27620 10192 27672 10198
rect 27620 10134 27672 10140
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 27436 9988 27488 9994
rect 27436 9930 27488 9936
rect 27528 9988 27580 9994
rect 27528 9930 27580 9936
rect 27344 9920 27396 9926
rect 27344 9862 27396 9868
rect 27356 7546 27384 9862
rect 27540 9518 27568 9930
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27436 9376 27488 9382
rect 27436 9318 27488 9324
rect 27448 8566 27476 9318
rect 27436 8560 27488 8566
rect 27436 8502 27488 8508
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 27632 6798 27660 9998
rect 27724 9625 27752 11018
rect 27710 9616 27766 9625
rect 27710 9551 27766 9560
rect 27724 9450 27752 9551
rect 27712 9444 27764 9450
rect 27712 9386 27764 9392
rect 27710 7576 27766 7585
rect 27710 7511 27766 7520
rect 27724 6905 27752 7511
rect 27816 7342 27844 14486
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 27908 13569 27936 14010
rect 28092 13734 28120 15592
rect 28172 15574 28224 15580
rect 28276 15026 28304 18702
rect 28448 17808 28500 17814
rect 28448 17750 28500 17756
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28368 14958 28396 17138
rect 28460 17105 28488 17750
rect 28446 17096 28502 17105
rect 28446 17031 28502 17040
rect 28460 15026 28488 17031
rect 28552 15638 28580 19246
rect 28736 17882 28764 21082
rect 28724 17876 28776 17882
rect 28724 17818 28776 17824
rect 28828 16561 28856 25094
rect 29516 25052 29824 25061
rect 29516 25050 29522 25052
rect 29578 25050 29602 25052
rect 29658 25050 29682 25052
rect 29738 25050 29762 25052
rect 29818 25050 29824 25052
rect 29578 24998 29580 25050
rect 29760 24998 29762 25050
rect 29516 24996 29522 24998
rect 29578 24996 29602 24998
rect 29658 24996 29682 24998
rect 29738 24996 29762 24998
rect 29818 24996 29824 24998
rect 29516 24987 29824 24996
rect 29516 23964 29824 23973
rect 29516 23962 29522 23964
rect 29578 23962 29602 23964
rect 29658 23962 29682 23964
rect 29738 23962 29762 23964
rect 29818 23962 29824 23964
rect 29578 23910 29580 23962
rect 29760 23910 29762 23962
rect 29516 23908 29522 23910
rect 29578 23908 29602 23910
rect 29658 23908 29682 23910
rect 29738 23908 29762 23910
rect 29818 23908 29824 23910
rect 29516 23899 29824 23908
rect 30208 23882 30236 25298
rect 30300 24818 30328 25842
rect 31128 25226 31156 26250
rect 31116 25220 31168 25226
rect 31116 25162 31168 25168
rect 30380 24948 30432 24954
rect 30380 24890 30432 24896
rect 30932 24948 30984 24954
rect 30932 24890 30984 24896
rect 30288 24812 30340 24818
rect 30288 24754 30340 24760
rect 30392 24682 30420 24890
rect 30380 24676 30432 24682
rect 30380 24618 30432 24624
rect 30208 23854 30328 23882
rect 30944 23866 30972 24890
rect 31024 24812 31076 24818
rect 31024 24754 31076 24760
rect 29276 23656 29328 23662
rect 29276 23598 29328 23604
rect 29000 22636 29052 22642
rect 29000 22578 29052 22584
rect 29012 20874 29040 22578
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 29000 20868 29052 20874
rect 29000 20810 29052 20816
rect 28908 20800 28960 20806
rect 28908 20742 28960 20748
rect 28920 20618 28948 20742
rect 28920 20590 29040 20618
rect 29012 17202 29040 20590
rect 29104 18329 29132 21830
rect 29090 18320 29146 18329
rect 29090 18255 29146 18264
rect 29092 17876 29144 17882
rect 29092 17818 29144 17824
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 28908 16584 28960 16590
rect 28814 16552 28870 16561
rect 28908 16526 28960 16532
rect 28814 16487 28870 16496
rect 28724 15904 28776 15910
rect 28724 15846 28776 15852
rect 28736 15706 28764 15846
rect 28724 15700 28776 15706
rect 28724 15642 28776 15648
rect 28540 15632 28592 15638
rect 28540 15574 28592 15580
rect 28828 15450 28856 16487
rect 28920 16454 28948 16526
rect 28908 16448 28960 16454
rect 28908 16390 28960 16396
rect 29000 16448 29052 16454
rect 29000 16390 29052 16396
rect 28906 16008 28962 16017
rect 29012 15994 29040 16390
rect 28962 15966 29040 15994
rect 28906 15943 28962 15952
rect 28920 15570 28948 15943
rect 28908 15564 28960 15570
rect 28908 15506 28960 15512
rect 28736 15422 28856 15450
rect 28906 15464 28962 15473
rect 28448 15020 28500 15026
rect 28448 14962 28500 14968
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28460 14822 28488 14962
rect 28448 14816 28500 14822
rect 28448 14758 28500 14764
rect 28448 14272 28500 14278
rect 28448 14214 28500 14220
rect 28460 14006 28488 14214
rect 28448 14000 28500 14006
rect 28448 13942 28500 13948
rect 28080 13728 28132 13734
rect 28080 13670 28132 13676
rect 27894 13560 27950 13569
rect 27894 13495 27950 13504
rect 27988 13388 28040 13394
rect 27988 13330 28040 13336
rect 28000 12918 28028 13330
rect 27988 12912 28040 12918
rect 27988 12854 28040 12860
rect 28092 12850 28120 13670
rect 28172 13252 28224 13258
rect 28172 13194 28224 13200
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 27896 12232 27948 12238
rect 27896 12174 27948 12180
rect 27908 11694 27936 12174
rect 28184 11830 28212 13194
rect 28448 13184 28500 13190
rect 28448 13126 28500 13132
rect 28356 12912 28408 12918
rect 28356 12854 28408 12860
rect 28264 12844 28316 12850
rect 28264 12786 28316 12792
rect 28172 11824 28224 11830
rect 28172 11766 28224 11772
rect 27896 11688 27948 11694
rect 27896 11630 27948 11636
rect 27908 11393 27936 11630
rect 28276 11506 28304 12786
rect 28368 12306 28396 12854
rect 28356 12300 28408 12306
rect 28356 12242 28408 12248
rect 28092 11478 28304 11506
rect 27894 11384 27950 11393
rect 27894 11319 27950 11328
rect 27908 11218 27936 11319
rect 27896 11212 27948 11218
rect 27896 11154 27948 11160
rect 27986 11112 28042 11121
rect 27986 11047 28042 11056
rect 27894 9752 27950 9761
rect 27894 9687 27950 9696
rect 27908 9654 27936 9687
rect 28000 9654 28028 11047
rect 28092 10470 28120 11478
rect 28264 11348 28316 11354
rect 28264 11290 28316 11296
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 28184 10742 28212 10950
rect 28172 10736 28224 10742
rect 28172 10678 28224 10684
rect 28276 10674 28304 11290
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 28080 10464 28132 10470
rect 28080 10406 28132 10412
rect 28092 9926 28120 10406
rect 28356 10056 28408 10062
rect 28356 9998 28408 10004
rect 28264 9988 28316 9994
rect 28264 9930 28316 9936
rect 28080 9920 28132 9926
rect 28132 9880 28212 9908
rect 28080 9862 28132 9868
rect 27896 9648 27948 9654
rect 27896 9590 27948 9596
rect 27988 9648 28040 9654
rect 27988 9590 28040 9596
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 27908 9217 27936 9454
rect 27894 9208 27950 9217
rect 27894 9143 27950 9152
rect 28078 8664 28134 8673
rect 28078 8599 28134 8608
rect 27896 8424 27948 8430
rect 27896 8366 27948 8372
rect 27986 8392 28042 8401
rect 27804 7336 27856 7342
rect 27804 7278 27856 7284
rect 27710 6896 27766 6905
rect 27908 6882 27936 8366
rect 27986 8327 28042 8336
rect 28000 7478 28028 8327
rect 28092 7993 28120 8599
rect 28184 8294 28212 9880
rect 28276 9761 28304 9930
rect 28262 9752 28318 9761
rect 28262 9687 28318 9696
rect 28368 9518 28396 9998
rect 28356 9512 28408 9518
rect 28356 9454 28408 9460
rect 28460 9364 28488 13126
rect 28552 11150 28580 14962
rect 28736 14906 28764 15422
rect 28906 15399 28962 15408
rect 28816 15360 28868 15366
rect 28816 15302 28868 15308
rect 28828 15026 28856 15302
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 28736 14878 28856 14906
rect 28724 14340 28776 14346
rect 28724 14282 28776 14288
rect 28736 14006 28764 14282
rect 28724 14000 28776 14006
rect 28724 13942 28776 13948
rect 28828 13308 28856 14878
rect 28920 14482 28948 15399
rect 29104 15026 29132 17818
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 29196 16250 29224 17070
rect 29184 16244 29236 16250
rect 29184 16186 29236 16192
rect 29182 15328 29238 15337
rect 29182 15263 29238 15272
rect 29092 15020 29144 15026
rect 29092 14962 29144 14968
rect 28908 14476 28960 14482
rect 28908 14418 28960 14424
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 29012 14278 29040 14418
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 28998 13696 29054 13705
rect 28920 13462 28948 13670
rect 28998 13631 29054 13640
rect 28908 13456 28960 13462
rect 28908 13398 28960 13404
rect 28828 13280 28948 13308
rect 28816 13184 28868 13190
rect 28816 13126 28868 13132
rect 28724 12844 28776 12850
rect 28724 12786 28776 12792
rect 28632 12300 28684 12306
rect 28632 12242 28684 12248
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28644 9738 28672 12242
rect 28736 12102 28764 12786
rect 28828 12782 28856 13126
rect 28816 12776 28868 12782
rect 28816 12718 28868 12724
rect 28920 12628 28948 13280
rect 28828 12600 28948 12628
rect 28724 12096 28776 12102
rect 28724 12038 28776 12044
rect 28828 11778 28856 12600
rect 29012 12442 29040 13631
rect 29090 13560 29146 13569
rect 29090 13495 29146 13504
rect 29104 12850 29132 13495
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 29000 12436 29052 12442
rect 29000 12378 29052 12384
rect 28908 12096 28960 12102
rect 28908 12038 28960 12044
rect 28920 11898 28948 12038
rect 29196 11898 29224 15263
rect 29288 14482 29316 23598
rect 29920 23316 29972 23322
rect 29920 23258 29972 23264
rect 29516 22876 29824 22885
rect 29516 22874 29522 22876
rect 29578 22874 29602 22876
rect 29658 22874 29682 22876
rect 29738 22874 29762 22876
rect 29818 22874 29824 22876
rect 29578 22822 29580 22874
rect 29760 22822 29762 22874
rect 29516 22820 29522 22822
rect 29578 22820 29602 22822
rect 29658 22820 29682 22822
rect 29738 22820 29762 22822
rect 29818 22820 29824 22822
rect 29516 22811 29824 22820
rect 29516 21788 29824 21797
rect 29516 21786 29522 21788
rect 29578 21786 29602 21788
rect 29658 21786 29682 21788
rect 29738 21786 29762 21788
rect 29818 21786 29824 21788
rect 29578 21734 29580 21786
rect 29760 21734 29762 21786
rect 29516 21732 29522 21734
rect 29578 21732 29602 21734
rect 29658 21732 29682 21734
rect 29738 21732 29762 21734
rect 29818 21732 29824 21734
rect 29516 21723 29824 21732
rect 29932 21570 29960 23258
rect 30012 22976 30064 22982
rect 30012 22918 30064 22924
rect 29840 21542 29960 21570
rect 29840 21146 29868 21542
rect 30024 21434 30052 22918
rect 30300 22166 30328 23854
rect 30932 23860 30984 23866
rect 30932 23802 30984 23808
rect 30472 23724 30524 23730
rect 30472 23666 30524 23672
rect 30380 23588 30432 23594
rect 30380 23530 30432 23536
rect 30288 22160 30340 22166
rect 30288 22102 30340 22108
rect 29932 21406 30052 21434
rect 29828 21140 29880 21146
rect 29828 21082 29880 21088
rect 29932 20806 29960 21406
rect 30012 21344 30064 21350
rect 30012 21286 30064 21292
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29920 20800 29972 20806
rect 29920 20742 29972 20748
rect 29380 17649 29408 20742
rect 29516 20700 29824 20709
rect 29516 20698 29522 20700
rect 29578 20698 29602 20700
rect 29658 20698 29682 20700
rect 29738 20698 29762 20700
rect 29818 20698 29824 20700
rect 29578 20646 29580 20698
rect 29760 20646 29762 20698
rect 29516 20644 29522 20646
rect 29578 20644 29602 20646
rect 29658 20644 29682 20646
rect 29738 20644 29762 20646
rect 29818 20644 29824 20646
rect 29516 20635 29824 20644
rect 30024 20534 30052 21286
rect 30196 21140 30248 21146
rect 30196 21082 30248 21088
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 30012 20528 30064 20534
rect 30012 20470 30064 20476
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 29516 19612 29824 19621
rect 29516 19610 29522 19612
rect 29578 19610 29602 19612
rect 29658 19610 29682 19612
rect 29738 19610 29762 19612
rect 29818 19610 29824 19612
rect 29578 19558 29580 19610
rect 29760 19558 29762 19610
rect 29516 19556 29522 19558
rect 29578 19556 29602 19558
rect 29658 19556 29682 19558
rect 29738 19556 29762 19558
rect 29818 19556 29824 19558
rect 29516 19547 29824 19556
rect 29516 18524 29824 18533
rect 29516 18522 29522 18524
rect 29578 18522 29602 18524
rect 29658 18522 29682 18524
rect 29738 18522 29762 18524
rect 29818 18522 29824 18524
rect 29578 18470 29580 18522
rect 29760 18470 29762 18522
rect 29516 18468 29522 18470
rect 29578 18468 29602 18470
rect 29658 18468 29682 18470
rect 29738 18468 29762 18470
rect 29818 18468 29824 18470
rect 29516 18459 29824 18468
rect 29366 17640 29422 17649
rect 29366 17575 29422 17584
rect 29516 17436 29824 17445
rect 29516 17434 29522 17436
rect 29578 17434 29602 17436
rect 29658 17434 29682 17436
rect 29738 17434 29762 17436
rect 29818 17434 29824 17436
rect 29578 17382 29580 17434
rect 29760 17382 29762 17434
rect 29516 17380 29522 17382
rect 29578 17380 29602 17382
rect 29658 17380 29682 17382
rect 29738 17380 29762 17382
rect 29818 17380 29824 17382
rect 29516 17371 29824 17380
rect 29734 17232 29790 17241
rect 29734 17167 29790 17176
rect 29748 17134 29776 17167
rect 29932 17134 29960 20334
rect 30116 19334 30144 20878
rect 30208 20097 30236 21082
rect 30300 20398 30328 22102
rect 30288 20392 30340 20398
rect 30288 20334 30340 20340
rect 30194 20088 30250 20097
rect 30194 20023 30250 20032
rect 30024 19306 30144 19334
rect 29736 17128 29788 17134
rect 29736 17070 29788 17076
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 29368 17060 29420 17066
rect 29368 17002 29420 17008
rect 29380 16046 29408 17002
rect 29920 16448 29972 16454
rect 29920 16390 29972 16396
rect 29516 16348 29824 16357
rect 29516 16346 29522 16348
rect 29578 16346 29602 16348
rect 29658 16346 29682 16348
rect 29738 16346 29762 16348
rect 29818 16346 29824 16348
rect 29578 16294 29580 16346
rect 29760 16294 29762 16346
rect 29516 16292 29522 16294
rect 29578 16292 29602 16294
rect 29658 16292 29682 16294
rect 29738 16292 29762 16294
rect 29818 16292 29824 16294
rect 29516 16283 29824 16292
rect 29932 16182 29960 16390
rect 29920 16176 29972 16182
rect 29920 16118 29972 16124
rect 29368 16040 29420 16046
rect 30024 15994 30052 19306
rect 30208 17898 30236 20023
rect 30208 17870 30328 17898
rect 30196 17672 30248 17678
rect 30196 17614 30248 17620
rect 30104 17196 30156 17202
rect 30104 17138 30156 17144
rect 30116 17105 30144 17138
rect 30102 17096 30158 17105
rect 30102 17031 30158 17040
rect 30104 16992 30156 16998
rect 30104 16934 30156 16940
rect 29368 15982 29420 15988
rect 29932 15966 30052 15994
rect 29932 15502 29960 15966
rect 29920 15496 29972 15502
rect 29920 15438 29972 15444
rect 29516 15260 29824 15269
rect 29516 15258 29522 15260
rect 29578 15258 29602 15260
rect 29658 15258 29682 15260
rect 29738 15258 29762 15260
rect 29818 15258 29824 15260
rect 29578 15206 29580 15258
rect 29760 15206 29762 15258
rect 29516 15204 29522 15206
rect 29578 15204 29602 15206
rect 29658 15204 29682 15206
rect 29738 15204 29762 15206
rect 29818 15204 29824 15206
rect 29516 15195 29824 15204
rect 29932 14958 29960 15438
rect 29920 14952 29972 14958
rect 29920 14894 29972 14900
rect 29276 14476 29328 14482
rect 29276 14418 29328 14424
rect 29920 14340 29972 14346
rect 29920 14282 29972 14288
rect 29276 14272 29328 14278
rect 29276 14214 29328 14220
rect 29288 12170 29316 14214
rect 29516 14172 29824 14181
rect 29516 14170 29522 14172
rect 29578 14170 29602 14172
rect 29658 14170 29682 14172
rect 29738 14170 29762 14172
rect 29818 14170 29824 14172
rect 29578 14118 29580 14170
rect 29760 14118 29762 14170
rect 29516 14116 29522 14118
rect 29578 14116 29602 14118
rect 29658 14116 29682 14118
rect 29738 14116 29762 14118
rect 29818 14116 29824 14118
rect 29516 14107 29824 14116
rect 29932 14074 29960 14282
rect 30012 14272 30064 14278
rect 30012 14214 30064 14220
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 29380 12850 29408 14010
rect 29920 13388 29972 13394
rect 29920 13330 29972 13336
rect 29516 13084 29824 13093
rect 29516 13082 29522 13084
rect 29578 13082 29602 13084
rect 29658 13082 29682 13084
rect 29738 13082 29762 13084
rect 29818 13082 29824 13084
rect 29578 13030 29580 13082
rect 29760 13030 29762 13082
rect 29516 13028 29522 13030
rect 29578 13028 29602 13030
rect 29658 13028 29682 13030
rect 29738 13028 29762 13030
rect 29818 13028 29824 13030
rect 29516 13019 29824 13028
rect 29932 12918 29960 13330
rect 30024 12918 30052 14214
rect 29920 12912 29972 12918
rect 29920 12854 29972 12860
rect 30012 12912 30064 12918
rect 30012 12854 30064 12860
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 29380 12306 29408 12786
rect 29368 12300 29420 12306
rect 29368 12242 29420 12248
rect 29276 12164 29328 12170
rect 29276 12106 29328 12112
rect 30012 12164 30064 12170
rect 30012 12106 30064 12112
rect 29920 12096 29972 12102
rect 29920 12038 29972 12044
rect 29516 11996 29824 12005
rect 29516 11994 29522 11996
rect 29578 11994 29602 11996
rect 29658 11994 29682 11996
rect 29738 11994 29762 11996
rect 29818 11994 29824 11996
rect 29578 11942 29580 11994
rect 29760 11942 29762 11994
rect 29516 11940 29522 11942
rect 29578 11940 29602 11942
rect 29658 11940 29682 11942
rect 29738 11940 29762 11942
rect 29818 11940 29824 11942
rect 29516 11931 29824 11940
rect 28908 11892 28960 11898
rect 28908 11834 28960 11840
rect 29184 11892 29236 11898
rect 29184 11834 29236 11840
rect 29460 11824 29512 11830
rect 28828 11750 28948 11778
rect 29460 11766 29512 11772
rect 28724 11620 28776 11626
rect 28724 11562 28776 11568
rect 28736 11529 28764 11562
rect 28722 11520 28778 11529
rect 28722 11455 28778 11464
rect 28816 11280 28868 11286
rect 28816 11222 28868 11228
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 28276 9336 28488 9364
rect 28552 9710 28672 9738
rect 28276 9194 28304 9336
rect 28552 9194 28580 9710
rect 28736 9625 28764 11086
rect 28828 9636 28856 11222
rect 28920 10064 28948 11750
rect 29092 11688 29144 11694
rect 29092 11630 29144 11636
rect 29104 10690 29132 11630
rect 29368 11552 29420 11558
rect 29368 11494 29420 11500
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 29184 11076 29236 11082
rect 29184 11018 29236 11024
rect 29017 10662 29132 10690
rect 29017 10656 29045 10662
rect 29012 10628 29045 10656
rect 28908 10058 28960 10064
rect 28908 10000 28960 10006
rect 29012 9704 29040 10628
rect 29092 10600 29144 10606
rect 29090 10568 29092 10577
rect 29144 10568 29146 10577
rect 29090 10503 29146 10512
rect 29196 9738 29224 11018
rect 29288 10810 29316 11290
rect 29276 10804 29328 10810
rect 29276 10746 29328 10752
rect 29380 10656 29408 11494
rect 29472 11354 29500 11766
rect 29644 11552 29696 11558
rect 29644 11494 29696 11500
rect 29460 11348 29512 11354
rect 29460 11290 29512 11296
rect 29656 11082 29684 11494
rect 29644 11076 29696 11082
rect 29644 11018 29696 11024
rect 29516 10908 29824 10917
rect 29516 10906 29522 10908
rect 29578 10906 29602 10908
rect 29658 10906 29682 10908
rect 29738 10906 29762 10908
rect 29818 10906 29824 10908
rect 29578 10854 29580 10906
rect 29760 10854 29762 10906
rect 29516 10852 29522 10854
rect 29578 10852 29602 10854
rect 29658 10852 29682 10854
rect 29738 10852 29762 10854
rect 29818 10852 29824 10854
rect 29516 10843 29824 10852
rect 29552 10736 29604 10742
rect 29552 10678 29604 10684
rect 29380 10628 29500 10656
rect 29472 10588 29500 10628
rect 29564 10588 29592 10678
rect 29472 10560 29592 10588
rect 29826 10568 29882 10577
rect 29826 10503 29882 10512
rect 29736 10192 29788 10198
rect 29736 10134 29788 10140
rect 29748 9926 29776 10134
rect 29840 9926 29868 10503
rect 29736 9920 29788 9926
rect 29736 9862 29788 9868
rect 29828 9920 29880 9926
rect 29828 9862 29880 9868
rect 29516 9820 29824 9829
rect 29516 9818 29522 9820
rect 29578 9818 29602 9820
rect 29658 9818 29682 9820
rect 29738 9818 29762 9820
rect 29818 9818 29824 9820
rect 29578 9766 29580 9818
rect 29760 9766 29762 9818
rect 29516 9764 29522 9766
rect 29578 9764 29602 9766
rect 29658 9764 29682 9766
rect 29738 9764 29762 9766
rect 29818 9764 29824 9766
rect 29516 9755 29824 9764
rect 29092 9716 29144 9722
rect 29012 9676 29092 9704
rect 29196 9710 29316 9738
rect 29092 9658 29144 9664
rect 29184 9648 29236 9654
rect 28722 9616 28778 9625
rect 28828 9608 28864 9636
rect 28722 9551 28778 9560
rect 28836 9500 28864 9608
rect 28998 9616 29054 9625
rect 29054 9574 29132 9602
rect 29184 9590 29236 9596
rect 28998 9551 29054 9560
rect 28836 9472 28948 9500
rect 28276 9166 28396 9194
rect 28552 9166 28672 9194
rect 28368 8548 28396 9166
rect 28540 9036 28592 9042
rect 28540 8978 28592 8984
rect 28448 8560 28500 8566
rect 28368 8520 28448 8548
rect 28448 8502 28500 8508
rect 28184 8266 28304 8294
rect 28078 7984 28134 7993
rect 28078 7919 28134 7928
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 27988 7472 28040 7478
rect 27988 7414 28040 7420
rect 27908 6854 28120 6882
rect 27710 6831 27766 6840
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 27344 6724 27396 6730
rect 27344 6666 27396 6672
rect 27356 5302 27384 6666
rect 27540 6458 27568 6734
rect 27528 6452 27580 6458
rect 27528 6394 27580 6400
rect 27816 5953 27844 6734
rect 27896 6384 27948 6390
rect 27896 6326 27948 6332
rect 27802 5944 27858 5953
rect 27802 5879 27858 5888
rect 27816 5778 27844 5879
rect 27804 5772 27856 5778
rect 27804 5714 27856 5720
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27620 5704 27672 5710
rect 27620 5646 27672 5652
rect 27344 5296 27396 5302
rect 27448 5273 27476 5646
rect 27528 5636 27580 5642
rect 27528 5578 27580 5584
rect 27344 5238 27396 5244
rect 27434 5264 27490 5273
rect 27540 5234 27568 5578
rect 27632 5545 27660 5646
rect 27804 5568 27856 5574
rect 27618 5536 27674 5545
rect 27618 5471 27674 5480
rect 27802 5536 27804 5545
rect 27856 5536 27858 5545
rect 27802 5471 27858 5480
rect 27434 5199 27490 5208
rect 27528 5228 27580 5234
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 27252 4684 27304 4690
rect 27252 4626 27304 4632
rect 27252 3936 27304 3942
rect 27252 3878 27304 3884
rect 27264 3534 27292 3878
rect 27356 3738 27384 4966
rect 27448 4826 27476 5199
rect 27528 5170 27580 5176
rect 27436 4820 27488 4826
rect 27436 4762 27488 4768
rect 27528 4480 27580 4486
rect 27528 4422 27580 4428
rect 27434 3768 27490 3777
rect 27344 3732 27396 3738
rect 27434 3703 27436 3712
rect 27344 3674 27396 3680
rect 27488 3703 27490 3712
rect 27436 3674 27488 3680
rect 27252 3528 27304 3534
rect 27252 3470 27304 3476
rect 27540 3466 27568 4422
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 27528 3460 27580 3466
rect 27528 3402 27580 3408
rect 27526 3224 27582 3233
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 27252 3188 27304 3194
rect 27526 3159 27582 3168
rect 27252 3130 27304 3136
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 27264 2310 27292 3130
rect 27540 3058 27568 3159
rect 27344 3052 27396 3058
rect 27528 3052 27580 3058
rect 27344 2994 27396 3000
rect 27448 3012 27528 3040
rect 27356 2310 27384 2994
rect 27448 2825 27476 3012
rect 27528 2994 27580 3000
rect 27620 2848 27672 2854
rect 27434 2816 27490 2825
rect 27434 2751 27490 2760
rect 27540 2796 27620 2802
rect 27540 2790 27672 2796
rect 27540 2774 27660 2790
rect 27540 2514 27568 2774
rect 27528 2508 27580 2514
rect 27528 2450 27580 2456
rect 27724 2378 27752 3878
rect 27908 3126 27936 6326
rect 28000 5710 28028 6734
rect 28092 5710 28120 6854
rect 28184 6662 28212 7482
rect 28276 6934 28304 8266
rect 28552 8242 28580 8978
rect 28644 8294 28672 9166
rect 28920 8838 28948 9472
rect 28998 9480 29054 9489
rect 28998 9415 29054 9424
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 28906 8664 28962 8673
rect 29012 8634 29040 9415
rect 28906 8599 28908 8608
rect 28960 8599 28962 8608
rect 29000 8628 29052 8634
rect 28908 8570 28960 8576
rect 29000 8570 29052 8576
rect 28908 8492 28960 8498
rect 29104 8480 29132 9574
rect 29196 9450 29224 9590
rect 29184 9444 29236 9450
rect 29184 9386 29236 9392
rect 29288 9110 29316 9710
rect 29460 9716 29512 9722
rect 29460 9658 29512 9664
rect 29552 9716 29604 9722
rect 29552 9658 29604 9664
rect 29276 9104 29328 9110
rect 29276 9046 29328 9052
rect 29472 8922 29500 9658
rect 29564 8974 29592 9658
rect 29932 9042 29960 12038
rect 30024 11830 30052 12106
rect 30012 11824 30064 11830
rect 30012 11766 30064 11772
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 30024 10062 30052 11086
rect 30012 10056 30064 10062
rect 30012 9998 30064 10004
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 30024 9518 30052 9862
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 30024 9042 30052 9454
rect 29920 9036 29972 9042
rect 29920 8978 29972 8984
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 28908 8434 28960 8440
rect 29012 8452 29132 8480
rect 29380 8894 29500 8922
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29920 8900 29972 8906
rect 28816 8356 28868 8362
rect 28816 8298 28868 8304
rect 28644 8266 28764 8294
rect 28368 8214 28580 8242
rect 28368 7410 28396 8214
rect 28630 8120 28686 8129
rect 28630 8055 28686 8064
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 28264 6928 28316 6934
rect 28264 6870 28316 6876
rect 28276 6798 28304 6870
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 28172 6656 28224 6662
rect 28172 6598 28224 6604
rect 28264 6656 28316 6662
rect 28264 6598 28316 6604
rect 28276 5817 28304 6598
rect 28262 5808 28318 5817
rect 28262 5743 28318 5752
rect 27988 5704 28040 5710
rect 27988 5646 28040 5652
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 28184 5234 28212 5306
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 28080 5092 28132 5098
rect 28080 5034 28132 5040
rect 28092 4214 28120 5034
rect 28368 4622 28396 7346
rect 28538 5944 28594 5953
rect 28538 5879 28594 5888
rect 28552 5778 28580 5879
rect 28644 5817 28672 8055
rect 28736 7750 28764 8266
rect 28828 8129 28856 8298
rect 28814 8120 28870 8129
rect 28814 8055 28870 8064
rect 28816 7880 28868 7886
rect 28920 7868 28948 8434
rect 29012 8362 29040 8452
rect 29380 8378 29408 8894
rect 29920 8842 29972 8848
rect 29516 8732 29824 8741
rect 29516 8730 29522 8732
rect 29578 8730 29602 8732
rect 29658 8730 29682 8732
rect 29738 8730 29762 8732
rect 29818 8730 29824 8732
rect 29578 8678 29580 8730
rect 29760 8678 29762 8730
rect 29516 8676 29522 8678
rect 29578 8676 29602 8678
rect 29658 8676 29682 8678
rect 29738 8676 29762 8678
rect 29818 8676 29824 8678
rect 29516 8667 29824 8676
rect 29932 8634 29960 8842
rect 29828 8628 29880 8634
rect 29828 8570 29880 8576
rect 29920 8628 29972 8634
rect 29920 8570 29972 8576
rect 29380 8362 29592 8378
rect 29000 8356 29052 8362
rect 29000 8298 29052 8304
rect 29092 8356 29144 8362
rect 29380 8356 29604 8362
rect 29380 8350 29552 8356
rect 29092 8298 29144 8304
rect 29552 8298 29604 8304
rect 29104 8022 29132 8298
rect 29840 8129 29868 8570
rect 29366 8120 29422 8129
rect 29366 8055 29422 8064
rect 29826 8120 29882 8129
rect 29826 8055 29882 8064
rect 29092 8016 29144 8022
rect 29092 7958 29144 7964
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 28868 7840 28948 7868
rect 28816 7822 28868 7828
rect 28724 7744 28776 7750
rect 28724 7686 28776 7692
rect 28630 5808 28686 5817
rect 28540 5772 28592 5778
rect 28630 5743 28686 5752
rect 28540 5714 28592 5720
rect 28448 5704 28500 5710
rect 28446 5672 28448 5681
rect 28500 5672 28502 5681
rect 28446 5607 28502 5616
rect 28540 5636 28592 5642
rect 28540 5578 28592 5584
rect 28552 5302 28580 5578
rect 28736 5574 28764 7686
rect 28724 5568 28776 5574
rect 28644 5528 28724 5556
rect 28540 5296 28592 5302
rect 28446 5264 28502 5273
rect 28540 5238 28592 5244
rect 28446 5199 28502 5208
rect 28460 5148 28488 5199
rect 28460 5120 28580 5148
rect 28552 4622 28580 5120
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 28184 4282 28212 4558
rect 28264 4548 28316 4554
rect 28264 4490 28316 4496
rect 28448 4548 28500 4554
rect 28448 4490 28500 4496
rect 28172 4276 28224 4282
rect 28172 4218 28224 4224
rect 28080 4208 28132 4214
rect 28080 4150 28132 4156
rect 28276 4010 28304 4490
rect 28264 4004 28316 4010
rect 28264 3946 28316 3952
rect 28276 3398 28304 3946
rect 28356 3732 28408 3738
rect 28356 3674 28408 3680
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 27896 3120 27948 3126
rect 27896 3062 27948 3068
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 28092 2854 28120 2994
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 27252 2304 27304 2310
rect 27252 2246 27304 2252
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 28368 800 28396 3674
rect 28460 3466 28488 4490
rect 28644 4078 28672 5528
rect 28724 5510 28776 5516
rect 28828 4865 28856 7822
rect 28908 7744 28960 7750
rect 28906 7712 28908 7721
rect 28960 7712 28962 7721
rect 28906 7647 28962 7656
rect 29012 7478 29040 7890
rect 29092 7744 29144 7750
rect 29092 7686 29144 7692
rect 29000 7472 29052 7478
rect 29000 7414 29052 7420
rect 29000 6996 29052 7002
rect 29000 6938 29052 6944
rect 29012 4978 29040 6938
rect 29104 6118 29132 7686
rect 29380 7478 29408 8055
rect 30024 7954 30052 8978
rect 30012 7948 30064 7954
rect 30012 7890 30064 7896
rect 29516 7644 29824 7653
rect 29516 7642 29522 7644
rect 29578 7642 29602 7644
rect 29658 7642 29682 7644
rect 29738 7642 29762 7644
rect 29818 7642 29824 7644
rect 29578 7590 29580 7642
rect 29760 7590 29762 7642
rect 29516 7588 29522 7590
rect 29578 7588 29602 7590
rect 29658 7588 29682 7590
rect 29738 7588 29762 7590
rect 29818 7588 29824 7590
rect 29516 7579 29824 7588
rect 29918 7576 29974 7585
rect 29918 7511 29974 7520
rect 29368 7472 29420 7478
rect 29368 7414 29420 7420
rect 29932 7313 29960 7511
rect 29918 7304 29974 7313
rect 29918 7239 29974 7248
rect 30010 6896 30066 6905
rect 30010 6831 30066 6840
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29092 6112 29144 6118
rect 29092 6054 29144 6060
rect 29288 5642 29316 6734
rect 29920 6656 29972 6662
rect 29920 6598 29972 6604
rect 29516 6556 29824 6565
rect 29516 6554 29522 6556
rect 29578 6554 29602 6556
rect 29658 6554 29682 6556
rect 29738 6554 29762 6556
rect 29818 6554 29824 6556
rect 29578 6502 29580 6554
rect 29760 6502 29762 6554
rect 29516 6500 29522 6502
rect 29578 6500 29602 6502
rect 29658 6500 29682 6502
rect 29738 6500 29762 6502
rect 29818 6500 29824 6502
rect 29516 6491 29824 6500
rect 29932 6390 29960 6598
rect 30024 6497 30052 6831
rect 30116 6746 30144 16934
rect 30208 15570 30236 17614
rect 30300 17542 30328 17870
rect 30288 17536 30340 17542
rect 30288 17478 30340 17484
rect 30392 17202 30420 23530
rect 30484 18834 30512 23666
rect 31036 22030 31064 24754
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31036 21554 31064 21966
rect 31128 21570 31156 25162
rect 31760 24744 31812 24750
rect 31760 24686 31812 24692
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31312 22030 31340 23802
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31404 22409 31432 22578
rect 31390 22400 31446 22409
rect 31390 22335 31446 22344
rect 31484 22092 31536 22098
rect 31484 22034 31536 22040
rect 31300 22024 31352 22030
rect 31300 21966 31352 21972
rect 31392 21616 31444 21622
rect 31024 21548 31076 21554
rect 31128 21542 31340 21570
rect 31392 21558 31444 21564
rect 31024 21490 31076 21496
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30852 21078 30880 21286
rect 30840 21072 30892 21078
rect 30840 21014 30892 21020
rect 31036 20942 31064 21490
rect 31312 21486 31340 21542
rect 31300 21480 31352 21486
rect 31300 21422 31352 21428
rect 31024 20936 31076 20942
rect 31024 20878 31076 20884
rect 30932 20800 30984 20806
rect 30932 20742 30984 20748
rect 30654 19544 30710 19553
rect 30654 19479 30710 19488
rect 30668 19446 30696 19479
rect 30656 19440 30708 19446
rect 30656 19382 30708 19388
rect 30746 19408 30802 19417
rect 30746 19343 30748 19352
rect 30800 19343 30802 19352
rect 30840 19372 30892 19378
rect 30748 19314 30800 19320
rect 30840 19314 30892 19320
rect 30852 18986 30880 19314
rect 30576 18958 30880 18986
rect 30472 18828 30524 18834
rect 30472 18770 30524 18776
rect 30380 17196 30432 17202
rect 30380 17138 30432 17144
rect 30380 17060 30432 17066
rect 30380 17002 30432 17008
rect 30392 16697 30420 17002
rect 30378 16688 30434 16697
rect 30378 16623 30434 16632
rect 30484 16454 30512 18770
rect 30576 17814 30604 18958
rect 30656 18896 30708 18902
rect 30654 18864 30656 18873
rect 30708 18864 30710 18873
rect 30654 18799 30710 18808
rect 30654 18728 30710 18737
rect 30654 18663 30710 18672
rect 30840 18692 30892 18698
rect 30668 18426 30696 18663
rect 30840 18634 30892 18640
rect 30748 18624 30800 18630
rect 30748 18566 30800 18572
rect 30656 18420 30708 18426
rect 30656 18362 30708 18368
rect 30564 17808 30616 17814
rect 30564 17750 30616 17756
rect 30576 17678 30604 17750
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30656 17604 30708 17610
rect 30656 17546 30708 17552
rect 30564 17196 30616 17202
rect 30564 17138 30616 17144
rect 30472 16448 30524 16454
rect 30472 16390 30524 16396
rect 30288 15904 30340 15910
rect 30288 15846 30340 15852
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 30208 14414 30236 15506
rect 30300 14958 30328 15846
rect 30484 15473 30512 16390
rect 30470 15464 30526 15473
rect 30470 15399 30526 15408
rect 30288 14952 30340 14958
rect 30288 14894 30340 14900
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 30196 14408 30248 14414
rect 30196 14350 30248 14356
rect 30208 13938 30236 14350
rect 30380 14068 30432 14074
rect 30380 14010 30432 14016
rect 30196 13932 30248 13938
rect 30196 13874 30248 13880
rect 30288 13456 30340 13462
rect 30288 13398 30340 13404
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30208 11150 30236 13262
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 30300 11098 30328 13398
rect 30392 12102 30420 14010
rect 30484 13190 30512 14418
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 30378 11928 30434 11937
rect 30378 11863 30434 11872
rect 30392 11218 30420 11863
rect 30380 11212 30432 11218
rect 30380 11154 30432 11160
rect 30300 11070 30420 11098
rect 30286 10976 30342 10985
rect 30286 10911 30342 10920
rect 30196 10464 30248 10470
rect 30196 10406 30248 10412
rect 30208 9926 30236 10406
rect 30196 9920 30248 9926
rect 30196 9862 30248 9868
rect 30194 9752 30250 9761
rect 30300 9722 30328 10911
rect 30194 9687 30250 9696
rect 30288 9716 30340 9722
rect 30208 9110 30236 9687
rect 30288 9658 30340 9664
rect 30286 9208 30342 9217
rect 30286 9143 30342 9152
rect 30196 9104 30248 9110
rect 30196 9046 30248 9052
rect 30300 8974 30328 9143
rect 30288 8968 30340 8974
rect 30288 8910 30340 8916
rect 30196 8900 30248 8906
rect 30196 8842 30248 8848
rect 30208 8566 30236 8842
rect 30286 8664 30342 8673
rect 30286 8599 30342 8608
rect 30196 8560 30248 8566
rect 30196 8502 30248 8508
rect 30300 8430 30328 8599
rect 30288 8424 30340 8430
rect 30288 8366 30340 8372
rect 30196 8288 30248 8294
rect 30196 8230 30248 8236
rect 30208 8090 30236 8230
rect 30196 8084 30248 8090
rect 30196 8026 30248 8032
rect 30286 7984 30342 7993
rect 30286 7919 30342 7928
rect 30300 7342 30328 7919
rect 30288 7336 30340 7342
rect 30288 7278 30340 7284
rect 30288 7200 30340 7206
rect 30288 7142 30340 7148
rect 30300 6866 30328 7142
rect 30288 6860 30340 6866
rect 30288 6802 30340 6808
rect 30116 6718 30236 6746
rect 30010 6488 30066 6497
rect 30010 6423 30066 6432
rect 29920 6384 29972 6390
rect 29920 6326 29972 6332
rect 29368 6248 29420 6254
rect 29368 6190 29420 6196
rect 29276 5636 29328 5642
rect 29276 5578 29328 5584
rect 29092 5568 29144 5574
rect 29092 5510 29144 5516
rect 29184 5568 29236 5574
rect 29184 5510 29236 5516
rect 29274 5536 29330 5545
rect 28920 4950 29040 4978
rect 28814 4856 28870 4865
rect 28814 4791 28870 4800
rect 28920 4570 28948 4950
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 29012 4690 29040 4762
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 28920 4542 29040 4570
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28632 4072 28684 4078
rect 28552 4032 28632 4060
rect 28448 3460 28500 3466
rect 28448 3402 28500 3408
rect 28552 2990 28580 4032
rect 28632 4014 28684 4020
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 28736 2650 28764 4082
rect 29012 3738 29040 4542
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 29000 3732 29052 3738
rect 29000 3674 29052 3680
rect 28920 3534 28948 3674
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 29104 3210 29132 5510
rect 29196 5166 29224 5510
rect 29274 5471 29330 5480
rect 29184 5160 29236 5166
rect 29184 5102 29236 5108
rect 29012 3182 29132 3210
rect 29012 3126 29040 3182
rect 29000 3120 29052 3126
rect 29000 3062 29052 3068
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 28920 1154 28948 2926
rect 29288 2310 29316 5471
rect 29380 5370 29408 6190
rect 30104 6112 30156 6118
rect 30104 6054 30156 6060
rect 30116 5846 30144 6054
rect 30012 5840 30064 5846
rect 30012 5782 30064 5788
rect 30104 5840 30156 5846
rect 30104 5782 30156 5788
rect 29920 5772 29972 5778
rect 29920 5714 29972 5720
rect 29516 5468 29824 5477
rect 29516 5466 29522 5468
rect 29578 5466 29602 5468
rect 29658 5466 29682 5468
rect 29738 5466 29762 5468
rect 29818 5466 29824 5468
rect 29578 5414 29580 5466
rect 29760 5414 29762 5466
rect 29516 5412 29522 5414
rect 29578 5412 29602 5414
rect 29658 5412 29682 5414
rect 29738 5412 29762 5414
rect 29818 5412 29824 5414
rect 29516 5403 29824 5412
rect 29932 5409 29960 5714
rect 29918 5400 29974 5409
rect 29368 5364 29420 5370
rect 29918 5335 29974 5344
rect 29368 5306 29420 5312
rect 29380 4622 29408 5306
rect 29920 5296 29972 5302
rect 29920 5238 29972 5244
rect 29368 4616 29420 4622
rect 29368 4558 29420 4564
rect 29380 4162 29408 4558
rect 29516 4380 29824 4389
rect 29516 4378 29522 4380
rect 29578 4378 29602 4380
rect 29658 4378 29682 4380
rect 29738 4378 29762 4380
rect 29818 4378 29824 4380
rect 29578 4326 29580 4378
rect 29760 4326 29762 4378
rect 29516 4324 29522 4326
rect 29578 4324 29602 4326
rect 29658 4324 29682 4326
rect 29738 4324 29762 4326
rect 29818 4324 29824 4326
rect 29516 4315 29824 4324
rect 29380 4134 29500 4162
rect 29472 4078 29500 4134
rect 29460 4072 29512 4078
rect 29460 4014 29512 4020
rect 29472 3602 29500 4014
rect 29932 3618 29960 5238
rect 30024 4690 30052 5782
rect 30104 5568 30156 5574
rect 30104 5510 30156 5516
rect 30116 5030 30144 5510
rect 30104 5024 30156 5030
rect 30104 4966 30156 4972
rect 30104 4820 30156 4826
rect 30104 4762 30156 4768
rect 30012 4684 30064 4690
rect 30012 4626 30064 4632
rect 30012 4548 30064 4554
rect 30012 4490 30064 4496
rect 30024 4214 30052 4490
rect 30012 4208 30064 4214
rect 30012 4150 30064 4156
rect 30010 4040 30066 4049
rect 30010 3975 30066 3984
rect 29460 3596 29512 3602
rect 29460 3538 29512 3544
rect 29656 3590 29960 3618
rect 29656 3534 29684 3590
rect 29644 3528 29696 3534
rect 29644 3470 29696 3476
rect 29516 3292 29824 3301
rect 29516 3290 29522 3292
rect 29578 3290 29602 3292
rect 29658 3290 29682 3292
rect 29738 3290 29762 3292
rect 29818 3290 29824 3292
rect 29578 3238 29580 3290
rect 29760 3238 29762 3290
rect 29516 3236 29522 3238
rect 29578 3236 29602 3238
rect 29658 3236 29682 3238
rect 29738 3236 29762 3238
rect 29818 3236 29824 3238
rect 29516 3227 29824 3236
rect 30024 3058 30052 3975
rect 30116 3534 30144 4762
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 30104 2848 30156 2854
rect 30104 2790 30156 2796
rect 30116 2446 30144 2790
rect 30208 2446 30236 6718
rect 30288 6452 30340 6458
rect 30288 6394 30340 6400
rect 30300 5370 30328 6394
rect 30392 5778 30420 11070
rect 30484 10538 30512 13126
rect 30576 12434 30604 17138
rect 30668 16658 30696 17546
rect 30656 16652 30708 16658
rect 30656 16594 30708 16600
rect 30668 15910 30696 16594
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30760 14346 30788 18566
rect 30852 18290 30880 18634
rect 30840 18284 30892 18290
rect 30840 18226 30892 18232
rect 30840 17196 30892 17202
rect 30840 17138 30892 17144
rect 30852 16590 30880 17138
rect 30840 16584 30892 16590
rect 30840 16526 30892 16532
rect 30944 16182 30972 20742
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 31036 18834 31064 19790
rect 31116 19372 31168 19378
rect 31116 19314 31168 19320
rect 31024 18828 31076 18834
rect 31024 18770 31076 18776
rect 31036 17746 31064 18770
rect 31024 17740 31076 17746
rect 31024 17682 31076 17688
rect 31036 17270 31064 17682
rect 31024 17264 31076 17270
rect 31024 17206 31076 17212
rect 30932 16176 30984 16182
rect 30932 16118 30984 16124
rect 30932 15972 30984 15978
rect 30932 15914 30984 15920
rect 30944 15706 30972 15914
rect 30932 15700 30984 15706
rect 30932 15642 30984 15648
rect 31128 15366 31156 19314
rect 31208 18692 31260 18698
rect 31208 18634 31260 18640
rect 31220 18222 31248 18634
rect 31312 18630 31340 21422
rect 31404 21010 31432 21558
rect 31496 21486 31524 22034
rect 31772 21690 31800 24686
rect 32036 24064 32088 24070
rect 32036 24006 32088 24012
rect 31852 23520 31904 23526
rect 31852 23462 31904 23468
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31484 21480 31536 21486
rect 31484 21422 31536 21428
rect 31392 21004 31444 21010
rect 31392 20946 31444 20952
rect 31300 18624 31352 18630
rect 31300 18566 31352 18572
rect 31208 18216 31260 18222
rect 31208 18158 31260 18164
rect 31300 18080 31352 18086
rect 31300 18022 31352 18028
rect 31312 17746 31340 18022
rect 31300 17740 31352 17746
rect 31300 17682 31352 17688
rect 31208 17536 31260 17542
rect 31208 17478 31260 17484
rect 31220 15706 31248 17478
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 31208 15700 31260 15706
rect 31208 15642 31260 15648
rect 31312 15638 31340 16050
rect 31300 15632 31352 15638
rect 31300 15574 31352 15580
rect 31404 15502 31432 20946
rect 31772 20942 31800 21626
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31772 20754 31800 20878
rect 31680 20726 31800 20754
rect 31680 19922 31708 20726
rect 31668 19916 31720 19922
rect 31668 19858 31720 19864
rect 31864 19786 31892 23462
rect 32048 19786 32076 24006
rect 32128 22976 32180 22982
rect 32128 22918 32180 22924
rect 32140 22506 32168 22918
rect 32416 22778 32444 26250
rect 32772 25696 32824 25702
rect 32772 25638 32824 25644
rect 32588 25220 32640 25226
rect 32588 25162 32640 25168
rect 32600 24206 32628 25162
rect 32588 24200 32640 24206
rect 32588 24142 32640 24148
rect 32404 22772 32456 22778
rect 32404 22714 32456 22720
rect 32128 22500 32180 22506
rect 32128 22442 32180 22448
rect 32600 22234 32628 24142
rect 32588 22228 32640 22234
rect 32588 22170 32640 22176
rect 32600 22094 32628 22170
rect 32784 22137 32812 25638
rect 33324 25424 33376 25430
rect 33324 25366 33376 25372
rect 32956 24132 33008 24138
rect 32956 24074 33008 24080
rect 32968 23662 32996 24074
rect 33048 23724 33100 23730
rect 33048 23666 33100 23672
rect 32956 23656 33008 23662
rect 32956 23598 33008 23604
rect 33060 23050 33088 23666
rect 33048 23044 33100 23050
rect 33048 22986 33100 22992
rect 32956 22636 33008 22642
rect 32956 22578 33008 22584
rect 32770 22128 32826 22137
rect 32600 22066 32720 22094
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 31852 19780 31904 19786
rect 31852 19722 31904 19728
rect 32036 19780 32088 19786
rect 32036 19722 32088 19728
rect 32600 18426 32628 20402
rect 32692 20398 32720 22066
rect 32770 22063 32826 22072
rect 32772 21888 32824 21894
rect 32864 21888 32916 21894
rect 32772 21830 32824 21836
rect 32862 21856 32864 21865
rect 32916 21856 32918 21865
rect 32784 20777 32812 21830
rect 32862 21791 32918 21800
rect 32864 20868 32916 20874
rect 32864 20810 32916 20816
rect 32770 20768 32826 20777
rect 32770 20703 32826 20712
rect 32680 20392 32732 20398
rect 32680 20334 32732 20340
rect 32588 18420 32640 18426
rect 32588 18362 32640 18368
rect 31576 18352 31628 18358
rect 31628 18312 31800 18340
rect 31576 18294 31628 18300
rect 31484 18284 31536 18290
rect 31484 18226 31536 18232
rect 31496 16153 31524 18226
rect 31666 17912 31722 17921
rect 31666 17847 31722 17856
rect 31680 17134 31708 17847
rect 31772 17746 31800 18312
rect 32496 17808 32548 17814
rect 32494 17776 32496 17785
rect 32548 17776 32550 17785
rect 31760 17740 31812 17746
rect 32494 17711 32550 17720
rect 31760 17682 31812 17688
rect 31576 17128 31628 17134
rect 31574 17096 31576 17105
rect 31668 17128 31720 17134
rect 31628 17096 31630 17105
rect 31668 17070 31720 17076
rect 31574 17031 31630 17040
rect 32312 16516 32364 16522
rect 32312 16458 32364 16464
rect 31482 16144 31538 16153
rect 31482 16079 31538 16088
rect 31496 15502 31524 16079
rect 31574 16008 31630 16017
rect 31574 15943 31630 15952
rect 31392 15496 31444 15502
rect 31392 15438 31444 15444
rect 31484 15496 31536 15502
rect 31484 15438 31536 15444
rect 31588 15434 31616 15943
rect 31760 15632 31812 15638
rect 31680 15592 31760 15620
rect 31576 15428 31628 15434
rect 31576 15370 31628 15376
rect 31116 15360 31168 15366
rect 31116 15302 31168 15308
rect 31680 15162 31708 15592
rect 31760 15574 31812 15580
rect 32220 15496 32272 15502
rect 32220 15438 32272 15444
rect 32036 15360 32088 15366
rect 32036 15302 32088 15308
rect 32128 15360 32180 15366
rect 32128 15302 32180 15308
rect 31668 15156 31720 15162
rect 31668 15098 31720 15104
rect 31392 15088 31444 15094
rect 31392 15030 31444 15036
rect 31024 14952 31076 14958
rect 31024 14894 31076 14900
rect 31036 14482 31064 14894
rect 31116 14816 31168 14822
rect 31116 14758 31168 14764
rect 31024 14476 31076 14482
rect 31024 14418 31076 14424
rect 30748 14340 30800 14346
rect 30748 14282 30800 14288
rect 30760 13138 30788 14282
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30852 13258 30880 14010
rect 31036 13410 31064 14418
rect 30944 13394 31064 13410
rect 30932 13388 31064 13394
rect 30984 13382 31064 13388
rect 30932 13330 30984 13336
rect 30840 13252 30892 13258
rect 30840 13194 30892 13200
rect 30760 13110 31064 13138
rect 30748 12640 30800 12646
rect 30748 12582 30800 12588
rect 30576 12406 30696 12434
rect 30564 12096 30616 12102
rect 30564 12038 30616 12044
rect 30576 11762 30604 12038
rect 30564 11756 30616 11762
rect 30564 11698 30616 11704
rect 30564 11552 30616 11558
rect 30564 11494 30616 11500
rect 30576 11014 30604 11494
rect 30564 11008 30616 11014
rect 30564 10950 30616 10956
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30472 10532 30524 10538
rect 30472 10474 30524 10480
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30484 6662 30512 8842
rect 30576 8401 30604 10610
rect 30562 8392 30618 8401
rect 30562 8327 30618 8336
rect 30562 7712 30618 7721
rect 30562 7647 30618 7656
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30470 6352 30526 6361
rect 30470 6287 30526 6296
rect 30380 5772 30432 5778
rect 30380 5714 30432 5720
rect 30378 5672 30434 5681
rect 30378 5607 30434 5616
rect 30392 5574 30420 5607
rect 30484 5574 30512 6287
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30472 5568 30524 5574
rect 30472 5510 30524 5516
rect 30288 5364 30340 5370
rect 30288 5306 30340 5312
rect 30392 5114 30420 5510
rect 30470 5264 30526 5273
rect 30576 5234 30604 7647
rect 30470 5199 30526 5208
rect 30564 5228 30616 5234
rect 30300 5086 30420 5114
rect 30300 4554 30328 5086
rect 30380 5024 30432 5030
rect 30380 4966 30432 4972
rect 30288 4548 30340 4554
rect 30288 4490 30340 4496
rect 30392 4078 30420 4966
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 30484 3466 30512 5199
rect 30564 5170 30616 5176
rect 30472 3460 30524 3466
rect 30472 3402 30524 3408
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30104 2440 30156 2446
rect 30104 2382 30156 2388
rect 30196 2440 30248 2446
rect 30196 2382 30248 2388
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29276 2304 29328 2310
rect 29276 2246 29328 2252
rect 29516 2204 29824 2213
rect 29516 2202 29522 2204
rect 29578 2202 29602 2204
rect 29658 2202 29682 2204
rect 29738 2202 29762 2204
rect 29818 2202 29824 2204
rect 29578 2150 29580 2202
rect 29760 2150 29762 2202
rect 29516 2148 29522 2150
rect 29578 2148 29602 2150
rect 29658 2148 29682 2150
rect 29738 2148 29762 2150
rect 29818 2148 29824 2150
rect 29516 2139 29824 2148
rect 29932 2106 29960 2314
rect 29920 2100 29972 2106
rect 29920 2042 29972 2048
rect 29736 2032 29788 2038
rect 29736 1974 29788 1980
rect 29748 1902 29776 1974
rect 29644 1896 29696 1902
rect 29644 1838 29696 1844
rect 29736 1896 29788 1902
rect 29736 1838 29788 1844
rect 29656 1698 29684 1838
rect 30392 1766 30420 2790
rect 30668 2650 30696 12406
rect 30760 11762 30788 12582
rect 31036 12434 31064 13110
rect 31128 12442 31156 14758
rect 31300 14340 31352 14346
rect 31300 14282 31352 14288
rect 30944 12406 31064 12434
rect 31116 12436 31168 12442
rect 30748 11756 30800 11762
rect 30748 11698 30800 11704
rect 30746 10840 30802 10849
rect 30746 10775 30802 10784
rect 30760 10305 30788 10775
rect 30746 10296 30802 10305
rect 30746 10231 30802 10240
rect 30760 10062 30788 10231
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 30838 9616 30894 9625
rect 30838 9551 30894 9560
rect 30748 9172 30800 9178
rect 30748 9114 30800 9120
rect 30760 8838 30788 9114
rect 30748 8832 30800 8838
rect 30748 8774 30800 8780
rect 30760 6866 30788 8774
rect 30748 6860 30800 6866
rect 30748 6802 30800 6808
rect 30748 5840 30800 5846
rect 30748 5782 30800 5788
rect 30760 4865 30788 5782
rect 30852 5234 30880 9551
rect 30944 7721 30972 12406
rect 31116 12378 31168 12384
rect 31128 11778 31156 12378
rect 31036 11750 31156 11778
rect 31036 11082 31064 11750
rect 31116 11688 31168 11694
rect 31208 11688 31260 11694
rect 31116 11630 31168 11636
rect 31206 11656 31208 11665
rect 31260 11656 31262 11665
rect 31024 11076 31076 11082
rect 31024 11018 31076 11024
rect 31024 10124 31076 10130
rect 31024 10066 31076 10072
rect 31036 9722 31064 10066
rect 31024 9716 31076 9722
rect 31024 9658 31076 9664
rect 31024 9512 31076 9518
rect 31024 9454 31076 9460
rect 31036 9178 31064 9454
rect 31024 9172 31076 9178
rect 31024 9114 31076 9120
rect 31022 9072 31078 9081
rect 31022 9007 31078 9016
rect 31036 8809 31064 9007
rect 31022 8800 31078 8809
rect 31022 8735 31078 8744
rect 31036 8566 31064 8735
rect 31024 8560 31076 8566
rect 31024 8502 31076 8508
rect 30930 7712 30986 7721
rect 30930 7647 30986 7656
rect 31024 7540 31076 7546
rect 31024 7482 31076 7488
rect 31036 7041 31064 7482
rect 31022 7032 31078 7041
rect 31022 6967 31078 6976
rect 30930 6896 30986 6905
rect 30930 6831 30986 6840
rect 30944 6730 30972 6831
rect 30932 6724 30984 6730
rect 30932 6666 30984 6672
rect 30932 5772 30984 5778
rect 30932 5714 30984 5720
rect 30840 5228 30892 5234
rect 30840 5170 30892 5176
rect 30746 4856 30802 4865
rect 30746 4791 30802 4800
rect 30852 3942 30880 5170
rect 30944 5166 30972 5714
rect 31022 5400 31078 5409
rect 31022 5335 31078 5344
rect 30932 5160 30984 5166
rect 30932 5102 30984 5108
rect 31036 4758 31064 5335
rect 31128 5273 31156 11630
rect 31206 11591 31262 11600
rect 31312 11354 31340 14282
rect 31404 12102 31432 15030
rect 31760 14816 31812 14822
rect 31760 14758 31812 14764
rect 31484 14272 31536 14278
rect 31484 14214 31536 14220
rect 31576 14272 31628 14278
rect 31576 14214 31628 14220
rect 31496 12986 31524 14214
rect 31484 12980 31536 12986
rect 31484 12922 31536 12928
rect 31496 12102 31524 12922
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31484 12096 31536 12102
rect 31484 12038 31536 12044
rect 31404 11762 31432 12038
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31208 11212 31260 11218
rect 31208 11154 31260 11160
rect 31220 11121 31248 11154
rect 31206 11112 31262 11121
rect 31588 11082 31616 14214
rect 31772 13138 31800 14758
rect 31852 13864 31904 13870
rect 31852 13806 31904 13812
rect 31864 13258 31892 13806
rect 31852 13252 31904 13258
rect 31852 13194 31904 13200
rect 32048 13138 32076 15302
rect 31772 13110 31892 13138
rect 31760 12980 31812 12986
rect 31760 12922 31812 12928
rect 31772 12782 31800 12922
rect 31760 12776 31812 12782
rect 31760 12718 31812 12724
rect 31758 12608 31814 12617
rect 31758 12543 31814 12552
rect 31668 12368 31720 12374
rect 31668 12310 31720 12316
rect 31206 11047 31262 11056
rect 31300 11076 31352 11082
rect 31300 11018 31352 11024
rect 31576 11076 31628 11082
rect 31576 11018 31628 11024
rect 31208 10532 31260 10538
rect 31208 10474 31260 10480
rect 31220 8430 31248 10474
rect 31208 8424 31260 8430
rect 31206 8392 31208 8401
rect 31260 8392 31262 8401
rect 31206 8327 31262 8336
rect 31312 8265 31340 11018
rect 31484 11008 31536 11014
rect 31484 10950 31536 10956
rect 31392 10668 31444 10674
rect 31392 10610 31444 10616
rect 31404 10470 31432 10610
rect 31392 10464 31444 10470
rect 31392 10406 31444 10412
rect 31392 9920 31444 9926
rect 31392 9862 31444 9868
rect 31404 9761 31432 9862
rect 31390 9752 31446 9761
rect 31390 9687 31446 9696
rect 31496 9466 31524 10950
rect 31680 10266 31708 12310
rect 31772 12306 31800 12543
rect 31760 12300 31812 12306
rect 31760 12242 31812 12248
rect 31760 11824 31812 11830
rect 31760 11766 31812 11772
rect 31772 11218 31800 11766
rect 31760 11212 31812 11218
rect 31760 11154 31812 11160
rect 31864 10674 31892 13110
rect 31956 13110 32076 13138
rect 31852 10668 31904 10674
rect 31852 10610 31904 10616
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 31956 10062 31984 13110
rect 32034 12336 32090 12345
rect 32034 12271 32090 12280
rect 32048 11286 32076 12271
rect 32140 11694 32168 15302
rect 32128 11688 32180 11694
rect 32128 11630 32180 11636
rect 32036 11280 32088 11286
rect 32036 11222 32088 11228
rect 32140 11132 32168 11630
rect 32048 11104 32168 11132
rect 32048 10130 32076 11104
rect 32128 11008 32180 11014
rect 32128 10950 32180 10956
rect 32140 10470 32168 10950
rect 32128 10464 32180 10470
rect 32128 10406 32180 10412
rect 32036 10124 32088 10130
rect 32036 10066 32088 10072
rect 31944 10056 31996 10062
rect 31944 9998 31996 10004
rect 31852 9920 31904 9926
rect 31852 9862 31904 9868
rect 31668 9716 31720 9722
rect 31668 9658 31720 9664
rect 31496 9438 31616 9466
rect 31484 9376 31536 9382
rect 31390 9344 31446 9353
rect 31484 9318 31536 9324
rect 31390 9279 31446 9288
rect 31404 9081 31432 9279
rect 31390 9072 31446 9081
rect 31390 9007 31446 9016
rect 31392 8560 31444 8566
rect 31392 8502 31444 8508
rect 31298 8256 31354 8265
rect 31298 8191 31354 8200
rect 31404 8106 31432 8502
rect 31220 8078 31432 8106
rect 31220 7342 31248 8078
rect 31392 8016 31444 8022
rect 31392 7958 31444 7964
rect 31300 7744 31352 7750
rect 31300 7686 31352 7692
rect 31208 7336 31260 7342
rect 31208 7278 31260 7284
rect 31206 7032 31262 7041
rect 31206 6967 31262 6976
rect 31220 5574 31248 6967
rect 31312 6866 31340 7686
rect 31404 7274 31432 7958
rect 31392 7268 31444 7274
rect 31392 7210 31444 7216
rect 31496 6934 31524 9318
rect 31588 7698 31616 9438
rect 31680 8566 31708 9658
rect 31864 9217 31892 9862
rect 31944 9580 31996 9586
rect 31944 9522 31996 9528
rect 31850 9208 31906 9217
rect 31850 9143 31906 9152
rect 31760 9036 31812 9042
rect 31760 8978 31812 8984
rect 31668 8560 31720 8566
rect 31668 8502 31720 8508
rect 31668 8288 31720 8294
rect 31668 8230 31720 8236
rect 31680 7818 31708 8230
rect 31772 7954 31800 8978
rect 31864 8634 31892 9143
rect 31852 8628 31904 8634
rect 31852 8570 31904 8576
rect 31760 7948 31812 7954
rect 31760 7890 31812 7896
rect 31668 7812 31720 7818
rect 31668 7754 31720 7760
rect 31588 7670 31708 7698
rect 31576 7336 31628 7342
rect 31576 7278 31628 7284
rect 31392 6928 31444 6934
rect 31392 6870 31444 6876
rect 31484 6928 31536 6934
rect 31484 6870 31536 6876
rect 31300 6860 31352 6866
rect 31300 6802 31352 6808
rect 31404 6474 31432 6870
rect 31496 6798 31524 6870
rect 31484 6792 31536 6798
rect 31484 6734 31536 6740
rect 31312 6446 31432 6474
rect 31312 6322 31340 6446
rect 31392 6384 31444 6390
rect 31392 6326 31444 6332
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 31312 5710 31340 6054
rect 31300 5704 31352 5710
rect 31300 5646 31352 5652
rect 31208 5568 31260 5574
rect 31208 5510 31260 5516
rect 31114 5264 31170 5273
rect 31114 5199 31170 5208
rect 31300 5228 31352 5234
rect 31300 5170 31352 5176
rect 31024 4752 31076 4758
rect 31024 4694 31076 4700
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 30656 2644 30708 2650
rect 30656 2586 30708 2592
rect 31312 2514 31340 5170
rect 31404 4049 31432 6326
rect 31390 4040 31446 4049
rect 31390 3975 31446 3984
rect 31496 3398 31524 6734
rect 31588 3913 31616 7278
rect 31680 7206 31708 7670
rect 31760 7404 31812 7410
rect 31760 7346 31812 7352
rect 31668 7200 31720 7206
rect 31668 7142 31720 7148
rect 31680 7002 31708 7142
rect 31668 6996 31720 7002
rect 31668 6938 31720 6944
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 31680 4593 31708 6734
rect 31772 6644 31800 7346
rect 31864 6798 31892 8570
rect 31852 6792 31904 6798
rect 31852 6734 31904 6740
rect 31772 6616 31892 6644
rect 31760 6452 31812 6458
rect 31760 6394 31812 6400
rect 31772 5710 31800 6394
rect 31760 5704 31812 5710
rect 31760 5646 31812 5652
rect 31864 5556 31892 6616
rect 31772 5528 31892 5556
rect 31666 4584 31722 4593
rect 31666 4519 31722 4528
rect 31574 3904 31630 3913
rect 31574 3839 31630 3848
rect 31484 3392 31536 3398
rect 31484 3334 31536 3340
rect 31772 2825 31800 5528
rect 31956 5114 31984 9522
rect 32048 6798 32076 10066
rect 32126 8800 32182 8809
rect 32126 8735 32182 8744
rect 32036 6792 32088 6798
rect 32036 6734 32088 6740
rect 32036 5772 32088 5778
rect 32036 5714 32088 5720
rect 31864 5086 31984 5114
rect 31864 3058 31892 5086
rect 31944 5024 31996 5030
rect 31944 4966 31996 4972
rect 31956 4622 31984 4966
rect 32048 4690 32076 5714
rect 32140 5370 32168 8735
rect 32128 5364 32180 5370
rect 32128 5306 32180 5312
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 32036 4684 32088 4690
rect 32036 4626 32088 4632
rect 31944 4616 31996 4622
rect 31944 4558 31996 4564
rect 31944 4276 31996 4282
rect 31944 4218 31996 4224
rect 31956 3670 31984 4218
rect 32048 4146 32076 4626
rect 32140 4486 32168 5170
rect 32128 4480 32180 4486
rect 32128 4422 32180 4428
rect 32232 4162 32260 15438
rect 32324 15026 32352 16458
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 32324 14550 32352 14962
rect 32312 14544 32364 14550
rect 32312 14486 32364 14492
rect 32404 13388 32456 13394
rect 32404 13330 32456 13336
rect 32312 12096 32364 12102
rect 32312 12038 32364 12044
rect 32324 11830 32352 12038
rect 32312 11824 32364 11830
rect 32312 11766 32364 11772
rect 32416 11762 32444 13330
rect 32404 11756 32456 11762
rect 32404 11698 32456 11704
rect 32404 11280 32456 11286
rect 32404 11222 32456 11228
rect 32312 10736 32364 10742
rect 32312 10678 32364 10684
rect 32324 8634 32352 10678
rect 32416 10266 32444 11222
rect 32404 10260 32456 10266
rect 32404 10202 32456 10208
rect 32404 10056 32456 10062
rect 32404 9998 32456 10004
rect 32312 8628 32364 8634
rect 32312 8570 32364 8576
rect 32416 7546 32444 9998
rect 32508 8634 32536 17711
rect 32772 17672 32824 17678
rect 32772 17614 32824 17620
rect 32588 17536 32640 17542
rect 32588 17478 32640 17484
rect 32600 17270 32628 17478
rect 32784 17338 32812 17614
rect 32772 17332 32824 17338
rect 32772 17274 32824 17280
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32680 17128 32732 17134
rect 32680 17070 32732 17076
rect 32692 16658 32720 17070
rect 32680 16652 32732 16658
rect 32680 16594 32732 16600
rect 32784 16454 32812 17274
rect 32876 16726 32904 20810
rect 32968 17338 32996 22578
rect 33060 20058 33088 22986
rect 33140 22568 33192 22574
rect 33140 22510 33192 22516
rect 33152 22166 33180 22510
rect 33140 22160 33192 22166
rect 33140 22102 33192 22108
rect 33048 20052 33100 20058
rect 33048 19994 33100 20000
rect 33140 19508 33192 19514
rect 33140 19450 33192 19456
rect 33152 18834 33180 19450
rect 33232 19440 33284 19446
rect 33232 19382 33284 19388
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 33140 17672 33192 17678
rect 33140 17614 33192 17620
rect 32956 17332 33008 17338
rect 32956 17274 33008 17280
rect 33152 17218 33180 17614
rect 33060 17190 33180 17218
rect 32864 16720 32916 16726
rect 32864 16662 32916 16668
rect 32956 16516 33008 16522
rect 32956 16458 33008 16464
rect 32772 16448 32824 16454
rect 32772 16390 32824 16396
rect 32968 16114 32996 16458
rect 33060 16182 33088 17190
rect 33138 17096 33194 17105
rect 33138 17031 33194 17040
rect 33048 16176 33100 16182
rect 33048 16118 33100 16124
rect 32956 16108 33008 16114
rect 32956 16050 33008 16056
rect 32588 15904 32640 15910
rect 32588 15846 32640 15852
rect 32600 15094 32628 15846
rect 32956 15632 33008 15638
rect 32956 15574 33008 15580
rect 32680 15156 32732 15162
rect 32680 15098 32732 15104
rect 32864 15156 32916 15162
rect 32864 15098 32916 15104
rect 32588 15088 32640 15094
rect 32588 15030 32640 15036
rect 32692 14958 32720 15098
rect 32588 14952 32640 14958
rect 32588 14894 32640 14900
rect 32680 14952 32732 14958
rect 32680 14894 32732 14900
rect 32600 12434 32628 14894
rect 32680 14068 32732 14074
rect 32680 14010 32732 14016
rect 32692 12918 32720 14010
rect 32772 13864 32824 13870
rect 32772 13806 32824 13812
rect 32784 13530 32812 13806
rect 32772 13524 32824 13530
rect 32772 13466 32824 13472
rect 32876 13297 32904 15098
rect 32862 13288 32918 13297
rect 32862 13223 32918 13232
rect 32864 13184 32916 13190
rect 32864 13126 32916 13132
rect 32876 12986 32904 13126
rect 32864 12980 32916 12986
rect 32864 12922 32916 12928
rect 32680 12912 32732 12918
rect 32680 12854 32732 12860
rect 32864 12776 32916 12782
rect 32864 12718 32916 12724
rect 32600 12406 32720 12434
rect 32588 12096 32640 12102
rect 32588 12038 32640 12044
rect 32600 11694 32628 12038
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32600 11286 32628 11630
rect 32588 11280 32640 11286
rect 32588 11222 32640 11228
rect 32588 11144 32640 11150
rect 32588 11086 32640 11092
rect 32600 10606 32628 11086
rect 32692 10810 32720 12406
rect 32876 12306 32904 12718
rect 32864 12300 32916 12306
rect 32864 12242 32916 12248
rect 32772 12164 32824 12170
rect 32772 12106 32824 12112
rect 32784 10962 32812 12106
rect 32864 12096 32916 12102
rect 32864 12038 32916 12044
rect 32876 11082 32904 12038
rect 32864 11076 32916 11082
rect 32864 11018 32916 11024
rect 32784 10934 32904 10962
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32588 10600 32640 10606
rect 32588 10542 32640 10548
rect 32600 10305 32628 10542
rect 32586 10296 32642 10305
rect 32586 10231 32642 10240
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 32588 9512 32640 9518
rect 32588 9454 32640 9460
rect 32600 9110 32628 9454
rect 32588 9104 32640 9110
rect 32588 9046 32640 9052
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32692 7546 32720 10202
rect 32876 10146 32904 10934
rect 32968 10266 32996 15574
rect 33152 14414 33180 17031
rect 33244 16590 33272 19382
rect 33232 16584 33284 16590
rect 33232 16526 33284 16532
rect 33232 16448 33284 16454
rect 33232 16390 33284 16396
rect 33244 15586 33272 16390
rect 33336 16182 33364 25366
rect 33414 17640 33470 17649
rect 33414 17575 33470 17584
rect 33324 16176 33376 16182
rect 33324 16118 33376 16124
rect 33244 15558 33364 15586
rect 33232 15496 33284 15502
rect 33232 15438 33284 15444
rect 33244 15366 33272 15438
rect 33232 15360 33284 15366
rect 33232 15302 33284 15308
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 33336 14090 33364 15558
rect 33428 15366 33456 17575
rect 33508 16584 33560 16590
rect 33508 16526 33560 16532
rect 33520 15502 33548 16526
rect 33508 15496 33560 15502
rect 33508 15438 33560 15444
rect 33416 15360 33468 15366
rect 33416 15302 33468 15308
rect 33508 14408 33560 14414
rect 33508 14350 33560 14356
rect 33336 14062 33456 14090
rect 33324 14000 33376 14006
rect 33324 13942 33376 13948
rect 33048 13932 33100 13938
rect 33048 13874 33100 13880
rect 33060 13734 33088 13874
rect 33140 13864 33192 13870
rect 33140 13806 33192 13812
rect 33048 13728 33100 13734
rect 33046 13696 33048 13705
rect 33100 13696 33102 13705
rect 33046 13631 33102 13640
rect 33048 13524 33100 13530
rect 33048 13466 33100 13472
rect 33060 12850 33088 13466
rect 33152 12986 33180 13806
rect 33140 12980 33192 12986
rect 33140 12922 33192 12928
rect 33336 12850 33364 13942
rect 33428 13546 33456 14062
rect 33520 13870 33548 14350
rect 33508 13864 33560 13870
rect 33508 13806 33560 13812
rect 33428 13518 33548 13546
rect 33416 12980 33468 12986
rect 33416 12922 33468 12928
rect 33048 12844 33100 12850
rect 33048 12786 33100 12792
rect 33324 12844 33376 12850
rect 33324 12786 33376 12792
rect 33138 12744 33194 12753
rect 33138 12679 33194 12688
rect 33048 12436 33100 12442
rect 33048 12378 33100 12384
rect 33060 12170 33088 12378
rect 33152 12374 33180 12679
rect 33324 12640 33376 12646
rect 33324 12582 33376 12588
rect 33230 12472 33286 12481
rect 33230 12407 33286 12416
rect 33140 12368 33192 12374
rect 33140 12310 33192 12316
rect 33048 12164 33100 12170
rect 33048 12106 33100 12112
rect 33140 12164 33192 12170
rect 33140 12106 33192 12112
rect 33048 11756 33100 11762
rect 33048 11698 33100 11704
rect 32956 10260 33008 10266
rect 32956 10202 33008 10208
rect 32876 10118 32996 10146
rect 32772 10056 32824 10062
rect 32772 9998 32824 10004
rect 32784 9042 32812 9998
rect 32864 9988 32916 9994
rect 32864 9930 32916 9936
rect 32876 9897 32904 9930
rect 32862 9888 32918 9897
rect 32862 9823 32918 9832
rect 32772 9036 32824 9042
rect 32772 8978 32824 8984
rect 32864 8628 32916 8634
rect 32864 8570 32916 8576
rect 32404 7540 32456 7546
rect 32404 7482 32456 7488
rect 32680 7540 32732 7546
rect 32680 7482 32732 7488
rect 32678 7440 32734 7449
rect 32678 7375 32680 7384
rect 32732 7375 32734 7384
rect 32680 7346 32732 7352
rect 32404 7336 32456 7342
rect 32404 7278 32456 7284
rect 32416 5846 32444 7278
rect 32692 6798 32720 7346
rect 32876 7041 32904 8570
rect 32968 8430 32996 10118
rect 33060 9722 33088 11698
rect 33152 11694 33180 12106
rect 33140 11688 33192 11694
rect 33140 11630 33192 11636
rect 33152 11529 33180 11630
rect 33138 11520 33194 11529
rect 33138 11455 33194 11464
rect 33244 10554 33272 12407
rect 33336 11626 33364 12582
rect 33428 12306 33456 12922
rect 33416 12300 33468 12306
rect 33416 12242 33468 12248
rect 33416 11892 33468 11898
rect 33416 11834 33468 11840
rect 33324 11620 33376 11626
rect 33324 11562 33376 11568
rect 33322 11520 33378 11529
rect 33322 11455 33378 11464
rect 33152 10526 33272 10554
rect 33048 9716 33100 9722
rect 33048 9658 33100 9664
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 33046 8392 33102 8401
rect 33046 8327 33102 8336
rect 33060 8294 33088 8327
rect 33048 8288 33100 8294
rect 32954 8256 33010 8265
rect 33048 8230 33100 8236
rect 32954 8191 33010 8200
rect 32968 7818 32996 8191
rect 32956 7812 33008 7818
rect 32956 7754 33008 7760
rect 32862 7032 32918 7041
rect 32862 6967 32918 6976
rect 32680 6792 32732 6798
rect 32680 6734 32732 6740
rect 32772 6724 32824 6730
rect 32772 6666 32824 6672
rect 32678 6488 32734 6497
rect 32678 6423 32734 6432
rect 32692 6390 32720 6423
rect 32680 6384 32732 6390
rect 32600 6344 32680 6372
rect 32496 6316 32548 6322
rect 32496 6258 32548 6264
rect 32404 5840 32456 5846
rect 32404 5782 32456 5788
rect 32404 5228 32456 5234
rect 32404 5170 32456 5176
rect 32416 5001 32444 5170
rect 32402 4992 32458 5001
rect 32402 4927 32458 4936
rect 32036 4140 32088 4146
rect 32232 4134 32352 4162
rect 32036 4082 32088 4088
rect 31944 3664 31996 3670
rect 31944 3606 31996 3612
rect 32048 3602 32076 4082
rect 32128 4004 32180 4010
rect 32128 3946 32180 3952
rect 32036 3596 32088 3602
rect 32036 3538 32088 3544
rect 31852 3052 31904 3058
rect 31852 2994 31904 3000
rect 31758 2816 31814 2825
rect 31758 2751 31814 2760
rect 32048 2514 32076 3538
rect 32140 3194 32168 3946
rect 32128 3188 32180 3194
rect 32128 3130 32180 3136
rect 32324 2922 32352 4134
rect 32402 3904 32458 3913
rect 32402 3839 32458 3848
rect 32416 3602 32444 3839
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 32508 3126 32536 6258
rect 32600 6225 32628 6344
rect 32680 6326 32732 6332
rect 32680 6248 32732 6254
rect 32586 6216 32642 6225
rect 32680 6190 32732 6196
rect 32586 6151 32642 6160
rect 32692 6118 32720 6190
rect 32784 6118 32812 6666
rect 33060 6254 33088 8230
rect 33048 6248 33100 6254
rect 33048 6190 33100 6196
rect 32680 6112 32732 6118
rect 32680 6054 32732 6060
rect 32772 6112 32824 6118
rect 32772 6054 32824 6060
rect 32956 5636 33008 5642
rect 32956 5578 33008 5584
rect 32968 4078 32996 5578
rect 33048 5092 33100 5098
rect 33048 5034 33100 5040
rect 33060 4690 33088 5034
rect 33048 4684 33100 4690
rect 33048 4626 33100 4632
rect 32680 4072 32732 4078
rect 32680 4014 32732 4020
rect 32956 4072 33008 4078
rect 32956 4014 33008 4020
rect 32692 3913 32720 4014
rect 33152 3942 33180 10526
rect 33230 10296 33286 10305
rect 33230 10231 33286 10240
rect 33244 9518 33272 10231
rect 33336 9874 33364 11455
rect 33428 10062 33456 11834
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33336 9846 33456 9874
rect 33232 9512 33284 9518
rect 33232 9454 33284 9460
rect 33244 7954 33272 9454
rect 33324 9376 33376 9382
rect 33324 9318 33376 9324
rect 33336 9081 33364 9318
rect 33322 9072 33378 9081
rect 33322 9007 33378 9016
rect 33428 8634 33456 9846
rect 33416 8628 33468 8634
rect 33416 8570 33468 8576
rect 33324 8492 33376 8498
rect 33324 8434 33376 8440
rect 33336 8090 33364 8434
rect 33416 8356 33468 8362
rect 33416 8298 33468 8304
rect 33324 8084 33376 8090
rect 33324 8026 33376 8032
rect 33232 7948 33284 7954
rect 33232 7890 33284 7896
rect 33244 7410 33272 7890
rect 33232 7404 33284 7410
rect 33232 7346 33284 7352
rect 33322 5672 33378 5681
rect 33322 5607 33378 5616
rect 33140 3936 33192 3942
rect 32678 3904 32734 3913
rect 33140 3878 33192 3884
rect 32678 3839 32734 3848
rect 33048 3732 33100 3738
rect 33048 3674 33100 3680
rect 32496 3120 32548 3126
rect 32496 3062 32548 3068
rect 32312 2916 32364 2922
rect 32312 2858 32364 2864
rect 33060 2854 33088 3674
rect 33336 3398 33364 5607
rect 33428 5166 33456 8298
rect 33520 8129 33548 13518
rect 33612 10810 33640 26522
rect 34164 24818 34192 26726
rect 34277 26684 34585 26693
rect 34277 26682 34283 26684
rect 34339 26682 34363 26684
rect 34419 26682 34443 26684
rect 34499 26682 34523 26684
rect 34579 26682 34585 26684
rect 34339 26630 34341 26682
rect 34521 26630 34523 26682
rect 34277 26628 34283 26630
rect 34339 26628 34363 26630
rect 34419 26628 34443 26630
rect 34499 26628 34523 26630
rect 34579 26628 34585 26630
rect 34277 26619 34585 26628
rect 34624 26382 34652 28478
rect 36082 28478 36308 28506
rect 36082 28354 36138 28478
rect 34704 26512 34756 26518
rect 34704 26454 34756 26460
rect 35532 26512 35584 26518
rect 35532 26454 35584 26460
rect 34612 26376 34664 26382
rect 34612 26318 34664 26324
rect 34277 25596 34585 25605
rect 34277 25594 34283 25596
rect 34339 25594 34363 25596
rect 34419 25594 34443 25596
rect 34499 25594 34523 25596
rect 34579 25594 34585 25596
rect 34339 25542 34341 25594
rect 34521 25542 34523 25594
rect 34277 25540 34283 25542
rect 34339 25540 34363 25542
rect 34419 25540 34443 25542
rect 34499 25540 34523 25542
rect 34579 25540 34585 25542
rect 34277 25531 34585 25540
rect 34152 24812 34204 24818
rect 34152 24754 34204 24760
rect 34716 24750 34744 26454
rect 34888 25764 34940 25770
rect 34888 25706 34940 25712
rect 34900 24954 34928 25706
rect 34888 24948 34940 24954
rect 34888 24890 34940 24896
rect 34704 24744 34756 24750
rect 34704 24686 34756 24692
rect 34277 24508 34585 24517
rect 34277 24506 34283 24508
rect 34339 24506 34363 24508
rect 34419 24506 34443 24508
rect 34499 24506 34523 24508
rect 34579 24506 34585 24508
rect 34339 24454 34341 24506
rect 34521 24454 34523 24506
rect 34277 24452 34283 24454
rect 34339 24452 34363 24454
rect 34419 24452 34443 24454
rect 34499 24452 34523 24454
rect 34579 24452 34585 24454
rect 34277 24443 34585 24452
rect 34716 24410 34744 24686
rect 34704 24404 34756 24410
rect 34704 24346 34756 24352
rect 34716 23730 34744 24346
rect 34704 23724 34756 23730
rect 34704 23666 34756 23672
rect 34277 23420 34585 23429
rect 34277 23418 34283 23420
rect 34339 23418 34363 23420
rect 34419 23418 34443 23420
rect 34499 23418 34523 23420
rect 34579 23418 34585 23420
rect 34339 23366 34341 23418
rect 34521 23366 34523 23418
rect 34277 23364 34283 23366
rect 34339 23364 34363 23366
rect 34419 23364 34443 23366
rect 34499 23364 34523 23366
rect 34579 23364 34585 23366
rect 34277 23355 34585 23364
rect 33968 22500 34020 22506
rect 33968 22442 34020 22448
rect 33692 21004 33744 21010
rect 33692 20946 33744 20952
rect 33704 20534 33732 20946
rect 33692 20528 33744 20534
rect 33692 20470 33744 20476
rect 33704 19825 33732 20470
rect 33690 19816 33746 19825
rect 33690 19751 33746 19760
rect 33784 19440 33836 19446
rect 33784 19382 33836 19388
rect 33692 16448 33744 16454
rect 33692 16390 33744 16396
rect 33704 16250 33732 16390
rect 33692 16244 33744 16250
rect 33692 16186 33744 16192
rect 33690 16008 33746 16017
rect 33690 15943 33746 15952
rect 33704 14074 33732 15943
rect 33796 15570 33824 19382
rect 33980 18290 34008 22442
rect 34277 22332 34585 22341
rect 34277 22330 34283 22332
rect 34339 22330 34363 22332
rect 34419 22330 34443 22332
rect 34499 22330 34523 22332
rect 34579 22330 34585 22332
rect 34339 22278 34341 22330
rect 34521 22278 34523 22330
rect 34277 22276 34283 22278
rect 34339 22276 34363 22278
rect 34419 22276 34443 22278
rect 34499 22276 34523 22278
rect 34579 22276 34585 22278
rect 34277 22267 34585 22276
rect 34277 21244 34585 21253
rect 34277 21242 34283 21244
rect 34339 21242 34363 21244
rect 34419 21242 34443 21244
rect 34499 21242 34523 21244
rect 34579 21242 34585 21244
rect 34339 21190 34341 21242
rect 34521 21190 34523 21242
rect 34277 21188 34283 21190
rect 34339 21188 34363 21190
rect 34419 21188 34443 21190
rect 34499 21188 34523 21190
rect 34579 21188 34585 21190
rect 34277 21179 34585 21188
rect 34796 20392 34848 20398
rect 34796 20334 34848 20340
rect 34277 20156 34585 20165
rect 34277 20154 34283 20156
rect 34339 20154 34363 20156
rect 34419 20154 34443 20156
rect 34499 20154 34523 20156
rect 34579 20154 34585 20156
rect 34339 20102 34341 20154
rect 34521 20102 34523 20154
rect 34277 20100 34283 20102
rect 34339 20100 34363 20102
rect 34419 20100 34443 20102
rect 34499 20100 34523 20102
rect 34579 20100 34585 20102
rect 34277 20091 34585 20100
rect 34702 19408 34758 19417
rect 34702 19343 34758 19352
rect 34716 19174 34744 19343
rect 34612 19168 34664 19174
rect 34612 19110 34664 19116
rect 34704 19168 34756 19174
rect 34704 19110 34756 19116
rect 34277 19068 34585 19077
rect 34277 19066 34283 19068
rect 34339 19066 34363 19068
rect 34419 19066 34443 19068
rect 34499 19066 34523 19068
rect 34579 19066 34585 19068
rect 34339 19014 34341 19066
rect 34521 19014 34523 19066
rect 34277 19012 34283 19014
rect 34339 19012 34363 19014
rect 34419 19012 34443 19014
rect 34499 19012 34523 19014
rect 34579 19012 34585 19014
rect 34277 19003 34585 19012
rect 34060 18692 34112 18698
rect 34060 18634 34112 18640
rect 33968 18284 34020 18290
rect 33968 18226 34020 18232
rect 33968 17808 34020 17814
rect 33968 17750 34020 17756
rect 33980 17270 34008 17750
rect 33968 17264 34020 17270
rect 33968 17206 34020 17212
rect 33968 16584 34020 16590
rect 33968 16526 34020 16532
rect 33876 16448 33928 16454
rect 33876 16390 33928 16396
rect 33888 16046 33916 16390
rect 33876 16040 33928 16046
rect 33876 15982 33928 15988
rect 33784 15564 33836 15570
rect 33784 15506 33836 15512
rect 33692 14068 33744 14074
rect 33692 14010 33744 14016
rect 33692 13932 33744 13938
rect 33692 13874 33744 13880
rect 33704 13530 33732 13874
rect 33692 13524 33744 13530
rect 33692 13466 33744 13472
rect 33704 13326 33732 13466
rect 33692 13320 33744 13326
rect 33692 13262 33744 13268
rect 33796 12481 33824 15506
rect 33980 14958 34008 16526
rect 33968 14952 34020 14958
rect 33968 14894 34020 14900
rect 33980 14634 34008 14894
rect 33888 14606 34008 14634
rect 33888 13326 33916 14606
rect 33968 13932 34020 13938
rect 33968 13874 34020 13880
rect 33980 13569 34008 13874
rect 33966 13560 34022 13569
rect 33966 13495 34022 13504
rect 34072 13462 34100 18634
rect 34152 18216 34204 18222
rect 34152 18158 34204 18164
rect 34164 17354 34192 18158
rect 34277 17980 34585 17989
rect 34277 17978 34283 17980
rect 34339 17978 34363 17980
rect 34419 17978 34443 17980
rect 34499 17978 34523 17980
rect 34579 17978 34585 17980
rect 34339 17926 34341 17978
rect 34521 17926 34523 17978
rect 34277 17924 34283 17926
rect 34339 17924 34363 17926
rect 34419 17924 34443 17926
rect 34499 17924 34523 17926
rect 34579 17924 34585 17926
rect 34277 17915 34585 17924
rect 34624 17746 34652 19110
rect 34612 17740 34664 17746
rect 34612 17682 34664 17688
rect 34164 17326 34376 17354
rect 34348 17270 34376 17326
rect 34336 17264 34388 17270
rect 34150 17232 34206 17241
rect 34336 17206 34388 17212
rect 34150 17167 34152 17176
rect 34204 17167 34206 17176
rect 34152 17138 34204 17144
rect 34348 17134 34376 17206
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34277 16892 34585 16901
rect 34277 16890 34283 16892
rect 34339 16890 34363 16892
rect 34419 16890 34443 16892
rect 34499 16890 34523 16892
rect 34579 16890 34585 16892
rect 34339 16838 34341 16890
rect 34521 16838 34523 16890
rect 34277 16836 34283 16838
rect 34339 16836 34363 16838
rect 34419 16836 34443 16838
rect 34499 16836 34523 16838
rect 34579 16836 34585 16838
rect 34277 16827 34585 16836
rect 34336 16516 34388 16522
rect 34336 16458 34388 16464
rect 34152 16040 34204 16046
rect 34348 16017 34376 16458
rect 34704 16176 34756 16182
rect 34704 16118 34756 16124
rect 34152 15982 34204 15988
rect 34334 16008 34390 16017
rect 34164 15910 34192 15982
rect 34334 15943 34390 15952
rect 34152 15904 34204 15910
rect 34152 15846 34204 15852
rect 34164 15434 34192 15846
rect 34277 15804 34585 15813
rect 34277 15802 34283 15804
rect 34339 15802 34363 15804
rect 34419 15802 34443 15804
rect 34499 15802 34523 15804
rect 34579 15802 34585 15804
rect 34339 15750 34341 15802
rect 34521 15750 34523 15802
rect 34277 15748 34283 15750
rect 34339 15748 34363 15750
rect 34419 15748 34443 15750
rect 34499 15748 34523 15750
rect 34579 15748 34585 15750
rect 34277 15739 34585 15748
rect 34152 15428 34204 15434
rect 34152 15370 34204 15376
rect 34277 14716 34585 14725
rect 34277 14714 34283 14716
rect 34339 14714 34363 14716
rect 34419 14714 34443 14716
rect 34499 14714 34523 14716
rect 34579 14714 34585 14716
rect 34339 14662 34341 14714
rect 34521 14662 34523 14714
rect 34277 14660 34283 14662
rect 34339 14660 34363 14662
rect 34419 14660 34443 14662
rect 34499 14660 34523 14662
rect 34579 14660 34585 14662
rect 34277 14651 34585 14660
rect 34716 14074 34744 16118
rect 34808 15978 34836 20334
rect 34900 17202 34928 24890
rect 35256 24812 35308 24818
rect 35084 24772 35256 24800
rect 35084 24614 35112 24772
rect 35256 24754 35308 24760
rect 35072 24608 35124 24614
rect 35072 24550 35124 24556
rect 34980 24268 35032 24274
rect 34980 24210 35032 24216
rect 34992 23730 35020 24210
rect 35084 24206 35112 24550
rect 35072 24200 35124 24206
rect 35072 24142 35124 24148
rect 35084 23730 35112 24142
rect 35440 24064 35492 24070
rect 35440 24006 35492 24012
rect 34980 23724 35032 23730
rect 34980 23666 35032 23672
rect 35072 23724 35124 23730
rect 35072 23666 35124 23672
rect 35164 20868 35216 20874
rect 35164 20810 35216 20816
rect 35176 20602 35204 20810
rect 35164 20596 35216 20602
rect 35164 20538 35216 20544
rect 34980 19372 35032 19378
rect 34980 19314 35032 19320
rect 34888 17196 34940 17202
rect 34888 17138 34940 17144
rect 34886 16552 34942 16561
rect 34886 16487 34942 16496
rect 34796 15972 34848 15978
rect 34796 15914 34848 15920
rect 34900 15910 34928 16487
rect 34888 15904 34940 15910
rect 34888 15846 34940 15852
rect 34888 15020 34940 15026
rect 34888 14962 34940 14968
rect 34900 14550 34928 14962
rect 34888 14544 34940 14550
rect 34888 14486 34940 14492
rect 34612 14068 34664 14074
rect 34612 14010 34664 14016
rect 34704 14068 34756 14074
rect 34704 14010 34756 14016
rect 34244 14000 34296 14006
rect 34244 13942 34296 13948
rect 34256 13802 34284 13942
rect 34244 13796 34296 13802
rect 34244 13738 34296 13744
rect 34277 13628 34585 13637
rect 34277 13626 34283 13628
rect 34339 13626 34363 13628
rect 34419 13626 34443 13628
rect 34499 13626 34523 13628
rect 34579 13626 34585 13628
rect 34339 13574 34341 13626
rect 34521 13574 34523 13626
rect 34277 13572 34283 13574
rect 34339 13572 34363 13574
rect 34419 13572 34443 13574
rect 34499 13572 34523 13574
rect 34579 13572 34585 13574
rect 34277 13563 34585 13572
rect 33968 13456 34020 13462
rect 33968 13398 34020 13404
rect 34060 13456 34112 13462
rect 34060 13398 34112 13404
rect 33876 13320 33928 13326
rect 33876 13262 33928 13268
rect 33980 13274 34008 13398
rect 33980 13246 34100 13274
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 33876 12640 33928 12646
rect 33876 12582 33928 12588
rect 33782 12472 33838 12481
rect 33782 12407 33838 12416
rect 33692 12300 33744 12306
rect 33692 12242 33744 12248
rect 33600 10804 33652 10810
rect 33600 10746 33652 10752
rect 33704 10538 33732 12242
rect 33888 11082 33916 12582
rect 33980 11762 34008 12786
rect 33968 11756 34020 11762
rect 33968 11698 34020 11704
rect 33968 11552 34020 11558
rect 33968 11494 34020 11500
rect 33980 11121 34008 11494
rect 33966 11112 34022 11121
rect 33876 11076 33928 11082
rect 33966 11047 34022 11056
rect 33876 11018 33928 11024
rect 34072 10962 34100 13246
rect 34152 12640 34204 12646
rect 34150 12608 34152 12617
rect 34204 12608 34206 12617
rect 34150 12543 34206 12552
rect 34277 12540 34585 12549
rect 34277 12538 34283 12540
rect 34339 12538 34363 12540
rect 34419 12538 34443 12540
rect 34499 12538 34523 12540
rect 34579 12538 34585 12540
rect 34339 12486 34341 12538
rect 34521 12486 34523 12538
rect 34277 12484 34283 12486
rect 34339 12484 34363 12486
rect 34419 12484 34443 12486
rect 34499 12484 34523 12486
rect 34579 12484 34585 12486
rect 34277 12475 34585 12484
rect 34624 12238 34652 14010
rect 34900 13394 34928 14486
rect 34796 13388 34848 13394
rect 34796 13330 34848 13336
rect 34888 13388 34940 13394
rect 34888 13330 34940 13336
rect 34808 12764 34836 13330
rect 34888 12776 34940 12782
rect 34808 12736 34888 12764
rect 34888 12718 34940 12724
rect 34888 12640 34940 12646
rect 34888 12582 34940 12588
rect 34900 12442 34928 12582
rect 34888 12436 34940 12442
rect 34888 12378 34940 12384
rect 34992 12322 35020 19314
rect 35452 18970 35480 24006
rect 35440 18964 35492 18970
rect 35440 18906 35492 18912
rect 35164 17604 35216 17610
rect 35164 17546 35216 17552
rect 35072 16652 35124 16658
rect 35072 16594 35124 16600
rect 35084 16182 35112 16594
rect 35176 16522 35204 17546
rect 35256 17128 35308 17134
rect 35256 17070 35308 17076
rect 35268 16590 35296 17070
rect 35544 16674 35572 26454
rect 36280 26382 36308 28478
rect 37370 28478 37688 28506
rect 37370 28354 37426 28478
rect 37660 26586 37688 28478
rect 38948 28478 39358 28506
rect 37648 26580 37700 26586
rect 37648 26522 37700 26528
rect 36268 26376 36320 26382
rect 36268 26318 36320 26324
rect 37554 26344 37610 26353
rect 37554 26279 37556 26288
rect 37608 26279 37610 26288
rect 37556 26250 37608 26256
rect 37556 25900 37608 25906
rect 37556 25842 37608 25848
rect 36728 25492 36780 25498
rect 36728 25434 36780 25440
rect 36268 25288 36320 25294
rect 36268 25230 36320 25236
rect 36452 25288 36504 25294
rect 36452 25230 36504 25236
rect 36636 25288 36688 25294
rect 36636 25230 36688 25236
rect 36280 24818 36308 25230
rect 36268 24812 36320 24818
rect 36268 24754 36320 24760
rect 36464 24750 36492 25230
rect 36648 24818 36676 25230
rect 36740 24886 36768 25434
rect 36728 24880 36780 24886
rect 36728 24822 36780 24828
rect 36544 24812 36596 24818
rect 36544 24754 36596 24760
rect 36636 24812 36688 24818
rect 36636 24754 36688 24760
rect 35900 24744 35952 24750
rect 35900 24686 35952 24692
rect 36084 24744 36136 24750
rect 36084 24686 36136 24692
rect 36452 24744 36504 24750
rect 36452 24686 36504 24692
rect 35912 24274 35940 24686
rect 36096 24614 36124 24686
rect 36084 24608 36136 24614
rect 36084 24550 36136 24556
rect 36556 24290 36584 24754
rect 36648 24410 36676 24754
rect 36636 24404 36688 24410
rect 36636 24346 36688 24352
rect 35900 24268 35952 24274
rect 35900 24210 35952 24216
rect 36464 24262 36584 24290
rect 35912 23594 35940 24210
rect 36464 24206 36492 24262
rect 36740 24206 36768 24822
rect 36912 24744 36964 24750
rect 36912 24686 36964 24692
rect 36924 24206 36952 24686
rect 36452 24200 36504 24206
rect 36452 24142 36504 24148
rect 36728 24200 36780 24206
rect 36728 24142 36780 24148
rect 36912 24200 36964 24206
rect 36912 24142 36964 24148
rect 35900 23588 35952 23594
rect 35900 23530 35952 23536
rect 35624 23520 35676 23526
rect 35624 23462 35676 23468
rect 35636 22094 35664 23462
rect 36464 23338 36492 24142
rect 37096 24064 37148 24070
rect 37096 24006 37148 24012
rect 36464 23310 36584 23338
rect 35636 22066 35756 22094
rect 35624 19372 35676 19378
rect 35624 19314 35676 19320
rect 35636 18834 35664 19314
rect 35624 18828 35676 18834
rect 35624 18770 35676 18776
rect 35728 18766 35756 22066
rect 36084 21548 36136 21554
rect 36084 21490 36136 21496
rect 36096 20466 36124 21490
rect 36176 20868 36228 20874
rect 36176 20810 36228 20816
rect 36188 20602 36216 20810
rect 36176 20596 36228 20602
rect 36176 20538 36228 20544
rect 36084 20460 36136 20466
rect 36084 20402 36136 20408
rect 36452 19712 36504 19718
rect 36452 19654 36504 19660
rect 36464 19514 36492 19654
rect 36452 19508 36504 19514
rect 36452 19450 36504 19456
rect 35900 19440 35952 19446
rect 35900 19382 35952 19388
rect 35716 18760 35768 18766
rect 35716 18702 35768 18708
rect 35912 18222 35940 19382
rect 35900 18216 35952 18222
rect 35900 18158 35952 18164
rect 36452 18216 36504 18222
rect 36452 18158 36504 18164
rect 35900 17740 35952 17746
rect 35900 17682 35952 17688
rect 35716 17264 35768 17270
rect 35716 17206 35768 17212
rect 35544 16646 35664 16674
rect 35256 16584 35308 16590
rect 35256 16526 35308 16532
rect 35532 16584 35584 16590
rect 35532 16526 35584 16532
rect 35164 16516 35216 16522
rect 35164 16458 35216 16464
rect 35072 16176 35124 16182
rect 35072 16118 35124 16124
rect 35072 15564 35124 15570
rect 35072 15506 35124 15512
rect 35084 15094 35112 15506
rect 35072 15088 35124 15094
rect 35164 15088 35216 15094
rect 35072 15030 35124 15036
rect 35162 15056 35164 15065
rect 35216 15056 35218 15065
rect 35162 14991 35218 15000
rect 35268 14906 35296 16526
rect 35348 16244 35400 16250
rect 35348 16186 35400 16192
rect 35176 14878 35296 14906
rect 35176 13954 35204 14878
rect 35256 14340 35308 14346
rect 35256 14282 35308 14288
rect 35268 14074 35296 14282
rect 35256 14068 35308 14074
rect 35256 14010 35308 14016
rect 35072 13932 35124 13938
rect 35176 13926 35296 13954
rect 35072 13874 35124 13880
rect 35084 12442 35112 13874
rect 35268 12986 35296 13926
rect 35256 12980 35308 12986
rect 35256 12922 35308 12928
rect 35256 12844 35308 12850
rect 35256 12786 35308 12792
rect 35268 12646 35296 12786
rect 35256 12640 35308 12646
rect 35256 12582 35308 12588
rect 35072 12436 35124 12442
rect 35072 12378 35124 12384
rect 34900 12294 35020 12322
rect 35084 12306 35112 12378
rect 35072 12300 35124 12306
rect 34612 12232 34664 12238
rect 34612 12174 34664 12180
rect 34152 12164 34204 12170
rect 34152 12106 34204 12112
rect 34796 12164 34848 12170
rect 34796 12106 34848 12112
rect 34164 11286 34192 12106
rect 34808 11762 34836 12106
rect 34796 11756 34848 11762
rect 34716 11716 34796 11744
rect 34612 11688 34664 11694
rect 34612 11630 34664 11636
rect 34277 11452 34585 11461
rect 34277 11450 34283 11452
rect 34339 11450 34363 11452
rect 34419 11450 34443 11452
rect 34499 11450 34523 11452
rect 34579 11450 34585 11452
rect 34339 11398 34341 11450
rect 34521 11398 34523 11450
rect 34277 11396 34283 11398
rect 34339 11396 34363 11398
rect 34419 11396 34443 11398
rect 34499 11396 34523 11398
rect 34579 11396 34585 11398
rect 34277 11387 34585 11396
rect 34152 11280 34204 11286
rect 34152 11222 34204 11228
rect 34428 11076 34480 11082
rect 34428 11018 34480 11024
rect 33796 10934 34100 10962
rect 33692 10532 33744 10538
rect 33692 10474 33744 10480
rect 33600 10464 33652 10470
rect 33600 10406 33652 10412
rect 33612 8974 33640 10406
rect 33796 9654 33824 10934
rect 33876 10804 33928 10810
rect 33876 10746 33928 10752
rect 33784 9648 33836 9654
rect 33784 9590 33836 9596
rect 33690 9208 33746 9217
rect 33690 9143 33746 9152
rect 33704 8974 33732 9143
rect 33600 8968 33652 8974
rect 33600 8910 33652 8916
rect 33692 8968 33744 8974
rect 33692 8910 33744 8916
rect 33782 8936 33838 8945
rect 33612 8566 33640 8910
rect 33782 8871 33784 8880
rect 33836 8871 33838 8880
rect 33784 8842 33836 8848
rect 33888 8616 33916 10746
rect 34440 10742 34468 11018
rect 34428 10736 34480 10742
rect 34428 10678 34480 10684
rect 34520 10668 34572 10674
rect 34624 10656 34652 11630
rect 34572 10628 34652 10656
rect 34520 10610 34572 10616
rect 34152 10532 34204 10538
rect 34152 10474 34204 10480
rect 33966 10432 34022 10441
rect 33966 10367 34022 10376
rect 33980 10062 34008 10367
rect 34058 10296 34114 10305
rect 34058 10231 34114 10240
rect 34072 10130 34100 10231
rect 34060 10124 34112 10130
rect 34060 10066 34112 10072
rect 33968 10056 34020 10062
rect 33968 9998 34020 10004
rect 33968 9920 34020 9926
rect 33968 9862 34020 9868
rect 33704 8588 33916 8616
rect 33600 8560 33652 8566
rect 33600 8502 33652 8508
rect 33704 8242 33732 8588
rect 33876 8492 33928 8498
rect 33876 8434 33928 8440
rect 33612 8214 33732 8242
rect 33784 8288 33836 8294
rect 33784 8230 33836 8236
rect 33506 8120 33562 8129
rect 33506 8055 33562 8064
rect 33506 6896 33562 6905
rect 33506 6831 33562 6840
rect 33520 6730 33548 6831
rect 33508 6724 33560 6730
rect 33508 6666 33560 6672
rect 33520 5778 33548 6666
rect 33508 5772 33560 5778
rect 33508 5714 33560 5720
rect 33520 5302 33548 5714
rect 33612 5681 33640 8214
rect 33690 8120 33746 8129
rect 33690 8055 33746 8064
rect 33598 5672 33654 5681
rect 33598 5607 33654 5616
rect 33598 5536 33654 5545
rect 33598 5471 33654 5480
rect 33508 5296 33560 5302
rect 33508 5238 33560 5244
rect 33416 5160 33468 5166
rect 33416 5102 33468 5108
rect 33612 4214 33640 5471
rect 33600 4208 33652 4214
rect 33600 4150 33652 4156
rect 33324 3392 33376 3398
rect 33324 3334 33376 3340
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33416 3120 33468 3126
rect 33414 3088 33416 3097
rect 33468 3088 33470 3097
rect 33414 3023 33470 3032
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33048 2848 33100 2854
rect 33048 2790 33100 2796
rect 33140 2848 33192 2854
rect 33140 2790 33192 2796
rect 31300 2508 31352 2514
rect 31300 2450 31352 2456
rect 32036 2508 32088 2514
rect 32036 2450 32088 2456
rect 32588 2508 32640 2514
rect 32588 2450 32640 2456
rect 30748 2372 30800 2378
rect 30748 2314 30800 2320
rect 30380 1760 30432 1766
rect 30380 1702 30432 1708
rect 29644 1692 29696 1698
rect 29644 1634 29696 1640
rect 28908 1148 28960 1154
rect 28908 1090 28960 1096
rect 30760 950 30788 2314
rect 31668 2304 31720 2310
rect 31668 2246 31720 2252
rect 31680 1834 31708 2246
rect 32600 2038 32628 2450
rect 32588 2032 32640 2038
rect 32588 1974 32640 1980
rect 31668 1828 31720 1834
rect 31668 1770 31720 1776
rect 33152 950 33180 2790
rect 33230 2680 33286 2689
rect 33230 2615 33286 2624
rect 33244 2378 33272 2615
rect 33232 2372 33284 2378
rect 33232 2314 33284 2320
rect 33520 1902 33548 2926
rect 33508 1896 33560 1902
rect 33508 1838 33560 1844
rect 33612 1698 33640 3334
rect 33704 2650 33732 8055
rect 33796 4865 33824 8230
rect 33888 6390 33916 8434
rect 33980 7954 34008 9862
rect 34058 9616 34114 9625
rect 34058 9551 34114 9560
rect 34072 8838 34100 9551
rect 34060 8832 34112 8838
rect 34060 8774 34112 8780
rect 34060 8424 34112 8430
rect 34060 8366 34112 8372
rect 34072 8294 34100 8366
rect 34060 8288 34112 8294
rect 34060 8230 34112 8236
rect 34060 8084 34112 8090
rect 34060 8026 34112 8032
rect 33968 7948 34020 7954
rect 33968 7890 34020 7896
rect 34072 7478 34100 8026
rect 34164 8022 34192 10474
rect 34277 10364 34585 10373
rect 34277 10362 34283 10364
rect 34339 10362 34363 10364
rect 34419 10362 34443 10364
rect 34499 10362 34523 10364
rect 34579 10362 34585 10364
rect 34339 10310 34341 10362
rect 34521 10310 34523 10362
rect 34277 10308 34283 10310
rect 34339 10308 34363 10310
rect 34419 10308 34443 10310
rect 34499 10308 34523 10310
rect 34579 10308 34585 10310
rect 34277 10299 34585 10308
rect 34624 10130 34652 10628
rect 34612 10124 34664 10130
rect 34612 10066 34664 10072
rect 34716 9674 34744 11716
rect 34796 11698 34848 11704
rect 34796 10600 34848 10606
rect 34796 10542 34848 10548
rect 34520 9648 34572 9654
rect 34518 9616 34520 9625
rect 34624 9646 34744 9674
rect 34572 9616 34574 9625
rect 34518 9551 34574 9560
rect 34277 9276 34585 9285
rect 34277 9274 34283 9276
rect 34339 9274 34363 9276
rect 34419 9274 34443 9276
rect 34499 9274 34523 9276
rect 34579 9274 34585 9276
rect 34339 9222 34341 9274
rect 34521 9222 34523 9274
rect 34277 9220 34283 9222
rect 34339 9220 34363 9222
rect 34419 9220 34443 9222
rect 34499 9220 34523 9222
rect 34579 9220 34585 9222
rect 34277 9211 34585 9220
rect 34624 9110 34652 9646
rect 34704 9172 34756 9178
rect 34704 9114 34756 9120
rect 34612 9104 34664 9110
rect 34612 9046 34664 9052
rect 34610 8800 34666 8809
rect 34610 8735 34666 8744
rect 34277 8188 34585 8197
rect 34277 8186 34283 8188
rect 34339 8186 34363 8188
rect 34419 8186 34443 8188
rect 34499 8186 34523 8188
rect 34579 8186 34585 8188
rect 34339 8134 34341 8186
rect 34521 8134 34523 8186
rect 34277 8132 34283 8134
rect 34339 8132 34363 8134
rect 34419 8132 34443 8134
rect 34499 8132 34523 8134
rect 34579 8132 34585 8134
rect 34277 8123 34585 8132
rect 34520 8084 34572 8090
rect 34520 8026 34572 8032
rect 34152 8016 34204 8022
rect 34152 7958 34204 7964
rect 34532 7562 34560 8026
rect 34440 7534 34560 7562
rect 34060 7472 34112 7478
rect 34060 7414 34112 7420
rect 34440 7290 34468 7534
rect 34164 7262 34468 7290
rect 34060 6792 34112 6798
rect 34060 6734 34112 6740
rect 34072 6633 34100 6734
rect 34058 6624 34114 6633
rect 34058 6559 34114 6568
rect 33876 6384 33928 6390
rect 33876 6326 33928 6332
rect 33888 5166 33916 6326
rect 33968 6316 34020 6322
rect 33968 6258 34020 6264
rect 33980 5953 34008 6258
rect 33966 5944 34022 5953
rect 33966 5879 34022 5888
rect 33876 5160 33928 5166
rect 33876 5102 33928 5108
rect 33782 4856 33838 4865
rect 33782 4791 33838 4800
rect 33796 4554 33824 4791
rect 33784 4548 33836 4554
rect 33784 4490 33836 4496
rect 33980 3194 34008 5879
rect 34072 3534 34100 6559
rect 34164 6458 34192 7262
rect 34277 7100 34585 7109
rect 34277 7098 34283 7100
rect 34339 7098 34363 7100
rect 34419 7098 34443 7100
rect 34499 7098 34523 7100
rect 34579 7098 34585 7100
rect 34339 7046 34341 7098
rect 34521 7046 34523 7098
rect 34277 7044 34283 7046
rect 34339 7044 34363 7046
rect 34419 7044 34443 7046
rect 34499 7044 34523 7046
rect 34579 7044 34585 7046
rect 34277 7035 34585 7044
rect 34242 6896 34298 6905
rect 34242 6831 34298 6840
rect 34152 6452 34204 6458
rect 34152 6394 34204 6400
rect 34256 6254 34284 6831
rect 34244 6248 34296 6254
rect 34244 6190 34296 6196
rect 34152 6112 34204 6118
rect 34152 6054 34204 6060
rect 34164 5556 34192 6054
rect 34277 6012 34585 6021
rect 34277 6010 34283 6012
rect 34339 6010 34363 6012
rect 34419 6010 34443 6012
rect 34499 6010 34523 6012
rect 34579 6010 34585 6012
rect 34339 5958 34341 6010
rect 34521 5958 34523 6010
rect 34277 5956 34283 5958
rect 34339 5956 34363 5958
rect 34419 5956 34443 5958
rect 34499 5956 34523 5958
rect 34579 5956 34585 5958
rect 34277 5947 34585 5956
rect 34624 5710 34652 8735
rect 34716 8634 34744 9114
rect 34704 8628 34756 8634
rect 34704 8570 34756 8576
rect 34702 8120 34758 8129
rect 34702 8055 34758 8064
rect 34716 7886 34744 8055
rect 34704 7880 34756 7886
rect 34704 7822 34756 7828
rect 34704 7336 34756 7342
rect 34704 7278 34756 7284
rect 34716 6798 34744 7278
rect 34704 6792 34756 6798
rect 34704 6734 34756 6740
rect 34612 5704 34664 5710
rect 34612 5646 34664 5652
rect 34244 5568 34296 5574
rect 34164 5528 34244 5556
rect 34244 5510 34296 5516
rect 34808 5370 34836 10542
rect 34900 9042 34928 12294
rect 35072 12242 35124 12248
rect 35164 12164 35216 12170
rect 35164 12106 35216 12112
rect 34978 11792 35034 11801
rect 34978 11727 35034 11736
rect 34992 11354 35020 11727
rect 34980 11348 35032 11354
rect 34980 11290 35032 11296
rect 34980 10804 35032 10810
rect 34980 10746 35032 10752
rect 34888 9036 34940 9042
rect 34888 8978 34940 8984
rect 34888 8900 34940 8906
rect 34888 8842 34940 8848
rect 34900 8498 34928 8842
rect 34992 8673 35020 10746
rect 35176 10146 35204 12106
rect 35084 10118 35204 10146
rect 34978 8664 35034 8673
rect 34978 8599 35034 8608
rect 34888 8492 34940 8498
rect 34888 8434 34940 8440
rect 34888 8288 34940 8294
rect 34888 8230 34940 8236
rect 34900 6934 34928 8230
rect 34992 6984 35020 8599
rect 35084 7154 35112 10118
rect 35164 9988 35216 9994
rect 35164 9930 35216 9936
rect 35176 9178 35204 9930
rect 35360 9926 35388 16186
rect 35440 15904 35492 15910
rect 35440 15846 35492 15852
rect 35452 15609 35480 15846
rect 35438 15600 35494 15609
rect 35438 15535 35494 15544
rect 35440 12980 35492 12986
rect 35440 12922 35492 12928
rect 35348 9920 35400 9926
rect 35348 9862 35400 9868
rect 35254 9752 35310 9761
rect 35254 9687 35310 9696
rect 35164 9172 35216 9178
rect 35164 9114 35216 9120
rect 35164 9036 35216 9042
rect 35164 8978 35216 8984
rect 35176 8820 35204 8978
rect 35268 8974 35296 9687
rect 35360 9042 35388 9862
rect 35348 9036 35400 9042
rect 35348 8978 35400 8984
rect 35256 8968 35308 8974
rect 35256 8910 35308 8916
rect 35176 8792 35296 8820
rect 35164 8424 35216 8430
rect 35164 8366 35216 8372
rect 35176 8294 35204 8366
rect 35164 8288 35216 8294
rect 35164 8230 35216 8236
rect 35164 7948 35216 7954
rect 35164 7890 35216 7896
rect 35176 7585 35204 7890
rect 35268 7732 35296 8792
rect 35452 8566 35480 12922
rect 35544 10849 35572 16526
rect 35636 13734 35664 16646
rect 35728 13802 35756 17206
rect 35808 16108 35860 16114
rect 35808 16050 35860 16056
rect 35820 13852 35848 16050
rect 35912 15094 35940 17682
rect 36464 17066 36492 18158
rect 36452 17060 36504 17066
rect 36452 17002 36504 17008
rect 36360 16448 36412 16454
rect 36360 16390 36412 16396
rect 35992 15700 36044 15706
rect 35992 15642 36044 15648
rect 35900 15088 35952 15094
rect 35900 15030 35952 15036
rect 35900 13864 35952 13870
rect 35820 13824 35900 13852
rect 35900 13806 35952 13812
rect 35716 13796 35768 13802
rect 35716 13738 35768 13744
rect 35624 13728 35676 13734
rect 35624 13670 35676 13676
rect 35636 12918 35664 13670
rect 35624 12912 35676 12918
rect 35624 12854 35676 12860
rect 35530 10840 35586 10849
rect 35728 10810 35756 13738
rect 35912 13190 35940 13806
rect 35900 13184 35952 13190
rect 35900 13126 35952 13132
rect 36004 12442 36032 15642
rect 36372 14414 36400 16390
rect 36464 15638 36492 17002
rect 36452 15632 36504 15638
rect 36452 15574 36504 15580
rect 36360 14408 36412 14414
rect 36360 14350 36412 14356
rect 36452 13796 36504 13802
rect 36452 13738 36504 13744
rect 35992 12436 36044 12442
rect 36464 12434 36492 13738
rect 35992 12378 36044 12384
rect 36372 12406 36492 12434
rect 35900 12232 35952 12238
rect 35900 12174 35952 12180
rect 35912 11694 35940 12174
rect 36084 12096 36136 12102
rect 36084 12038 36136 12044
rect 35900 11688 35952 11694
rect 35900 11630 35952 11636
rect 36096 11354 36124 12038
rect 36084 11348 36136 11354
rect 36084 11290 36136 11296
rect 35992 11280 36044 11286
rect 35992 11222 36044 11228
rect 35530 10775 35586 10784
rect 35716 10804 35768 10810
rect 35716 10746 35768 10752
rect 35808 10464 35860 10470
rect 35728 10424 35808 10452
rect 35728 9897 35756 10424
rect 35808 10406 35860 10412
rect 35714 9888 35770 9897
rect 35714 9823 35770 9832
rect 35624 9580 35676 9586
rect 35624 9522 35676 9528
rect 35636 9110 35664 9522
rect 35624 9104 35676 9110
rect 35624 9046 35676 9052
rect 35532 9036 35584 9042
rect 35532 8978 35584 8984
rect 35440 8560 35492 8566
rect 35440 8502 35492 8508
rect 35348 8356 35400 8362
rect 35348 8298 35400 8304
rect 35360 7886 35388 8298
rect 35348 7880 35400 7886
rect 35348 7822 35400 7828
rect 35268 7704 35388 7732
rect 35162 7576 35218 7585
rect 35162 7511 35218 7520
rect 35256 7540 35308 7546
rect 35256 7482 35308 7488
rect 35084 7126 35204 7154
rect 34992 6956 35112 6984
rect 34888 6928 34940 6934
rect 34940 6888 35020 6916
rect 34888 6870 34940 6876
rect 34886 6760 34942 6769
rect 34886 6695 34942 6704
rect 34900 6662 34928 6695
rect 34888 6656 34940 6662
rect 34888 6598 34940 6604
rect 34888 6248 34940 6254
rect 34888 6190 34940 6196
rect 34900 5914 34928 6190
rect 34888 5908 34940 5914
rect 34888 5850 34940 5856
rect 34704 5364 34756 5370
rect 34704 5306 34756 5312
rect 34796 5364 34848 5370
rect 34796 5306 34848 5312
rect 34716 5030 34744 5306
rect 34704 5024 34756 5030
rect 34704 4966 34756 4972
rect 34277 4924 34585 4933
rect 34277 4922 34283 4924
rect 34339 4922 34363 4924
rect 34419 4922 34443 4924
rect 34499 4922 34523 4924
rect 34579 4922 34585 4924
rect 34339 4870 34341 4922
rect 34521 4870 34523 4922
rect 34277 4868 34283 4870
rect 34339 4868 34363 4870
rect 34419 4868 34443 4870
rect 34499 4868 34523 4870
rect 34579 4868 34585 4870
rect 34277 4859 34585 4868
rect 34428 4820 34480 4826
rect 34428 4762 34480 4768
rect 34440 4486 34468 4762
rect 34428 4480 34480 4486
rect 34428 4422 34480 4428
rect 34796 4480 34848 4486
rect 34796 4422 34848 4428
rect 34277 3836 34585 3845
rect 34277 3834 34283 3836
rect 34339 3834 34363 3836
rect 34419 3834 34443 3836
rect 34499 3834 34523 3836
rect 34579 3834 34585 3836
rect 34339 3782 34341 3834
rect 34521 3782 34523 3834
rect 34277 3780 34283 3782
rect 34339 3780 34363 3782
rect 34419 3780 34443 3782
rect 34499 3780 34523 3782
rect 34579 3780 34585 3782
rect 34277 3771 34585 3780
rect 34060 3528 34112 3534
rect 34060 3470 34112 3476
rect 33968 3188 34020 3194
rect 33968 3130 34020 3136
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 34072 2446 34100 3470
rect 34808 3466 34836 4422
rect 34992 4078 35020 6888
rect 35084 4622 35112 6956
rect 35072 4616 35124 4622
rect 35072 4558 35124 4564
rect 35176 4282 35204 7126
rect 35268 6769 35296 7482
rect 35254 6760 35310 6769
rect 35254 6695 35310 6704
rect 35256 6656 35308 6662
rect 35256 6598 35308 6604
rect 35268 6225 35296 6598
rect 35254 6216 35310 6225
rect 35254 6151 35310 6160
rect 35360 6100 35388 7704
rect 35268 6072 35388 6100
rect 35268 5234 35296 6072
rect 35348 5908 35400 5914
rect 35348 5850 35400 5856
rect 35256 5228 35308 5234
rect 35256 5170 35308 5176
rect 35360 4808 35388 5850
rect 35452 5710 35480 8502
rect 35544 8430 35572 8978
rect 35636 8974 35664 9046
rect 35624 8968 35676 8974
rect 35624 8910 35676 8916
rect 35624 8832 35676 8838
rect 35624 8774 35676 8780
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 35532 7744 35584 7750
rect 35532 7686 35584 7692
rect 35440 5704 35492 5710
rect 35440 5646 35492 5652
rect 35360 4780 35480 4808
rect 35452 4729 35480 4780
rect 35438 4720 35494 4729
rect 35438 4655 35494 4664
rect 35164 4276 35216 4282
rect 35164 4218 35216 4224
rect 35452 4214 35480 4655
rect 35440 4208 35492 4214
rect 35440 4150 35492 4156
rect 34980 4072 35032 4078
rect 34980 4014 35032 4020
rect 34888 3596 34940 3602
rect 34888 3538 34940 3544
rect 34796 3460 34848 3466
rect 34796 3402 34848 3408
rect 34704 3120 34756 3126
rect 34704 3062 34756 3068
rect 34150 2816 34206 2825
rect 34150 2751 34206 2760
rect 34060 2440 34112 2446
rect 34060 2382 34112 2388
rect 34072 2310 34100 2382
rect 34164 2378 34192 2751
rect 34277 2748 34585 2757
rect 34277 2746 34283 2748
rect 34339 2746 34363 2748
rect 34419 2746 34443 2748
rect 34499 2746 34523 2748
rect 34579 2746 34585 2748
rect 34339 2694 34341 2746
rect 34521 2694 34523 2746
rect 34277 2692 34283 2694
rect 34339 2692 34363 2694
rect 34419 2692 34443 2694
rect 34499 2692 34523 2694
rect 34579 2692 34585 2694
rect 34277 2683 34585 2692
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 34060 2304 34112 2310
rect 34060 2246 34112 2252
rect 33600 1692 33652 1698
rect 33600 1634 33652 1640
rect 34716 1329 34744 3062
rect 34900 3058 34928 3538
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 34702 1320 34758 1329
rect 34702 1255 34758 1264
rect 35176 1222 35204 3402
rect 35544 2582 35572 7686
rect 35636 6254 35664 8774
rect 35624 6248 35676 6254
rect 35624 6190 35676 6196
rect 35624 5568 35676 5574
rect 35624 5510 35676 5516
rect 35636 4214 35664 5510
rect 35728 5370 35756 9823
rect 35900 9036 35952 9042
rect 35900 8978 35952 8984
rect 35808 8016 35860 8022
rect 35808 7958 35860 7964
rect 35820 6798 35848 7958
rect 35912 7954 35940 8978
rect 36004 8498 36032 11222
rect 36268 11212 36320 11218
rect 36268 11154 36320 11160
rect 36174 10024 36230 10033
rect 36174 9959 36230 9968
rect 36188 9178 36216 9959
rect 36176 9172 36228 9178
rect 36176 9114 36228 9120
rect 35992 8492 36044 8498
rect 35992 8434 36044 8440
rect 35900 7948 35952 7954
rect 36280 7936 36308 11154
rect 35900 7890 35952 7896
rect 36096 7908 36308 7936
rect 36096 7562 36124 7908
rect 36266 7848 36322 7857
rect 36176 7812 36228 7818
rect 36266 7783 36268 7792
rect 36176 7754 36228 7760
rect 36320 7783 36322 7792
rect 36268 7754 36320 7760
rect 35912 7534 36124 7562
rect 36188 7546 36216 7754
rect 36176 7540 36228 7546
rect 35808 6792 35860 6798
rect 35808 6734 35860 6740
rect 35912 6497 35940 7534
rect 36176 7482 36228 7488
rect 35992 7472 36044 7478
rect 35992 7414 36044 7420
rect 36004 7002 36032 7414
rect 36082 7304 36138 7313
rect 36082 7239 36138 7248
rect 36096 7002 36124 7239
rect 35992 6996 36044 7002
rect 35992 6938 36044 6944
rect 36084 6996 36136 7002
rect 36084 6938 36136 6944
rect 35992 6792 36044 6798
rect 35992 6734 36044 6740
rect 36084 6792 36136 6798
rect 36084 6734 36136 6740
rect 35898 6488 35954 6497
rect 35898 6423 35954 6432
rect 35912 6202 35940 6423
rect 35820 6174 35940 6202
rect 36004 6186 36032 6734
rect 36096 6633 36124 6734
rect 36082 6624 36138 6633
rect 36082 6559 36138 6568
rect 36174 6352 36230 6361
rect 36174 6287 36176 6296
rect 36228 6287 36230 6296
rect 36176 6258 36228 6264
rect 35992 6180 36044 6186
rect 35716 5364 35768 5370
rect 35716 5306 35768 5312
rect 35716 5228 35768 5234
rect 35716 5170 35768 5176
rect 35624 4208 35676 4214
rect 35624 4150 35676 4156
rect 35532 2576 35584 2582
rect 35532 2518 35584 2524
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35164 1216 35216 1222
rect 35164 1158 35216 1164
rect 29644 944 29696 950
rect 29644 886 29696 892
rect 30748 944 30800 950
rect 30748 886 30800 892
rect 31576 944 31628 950
rect 31576 886 31628 892
rect 33140 944 33192 950
rect 33140 886 33192 892
rect 33508 944 33560 950
rect 33508 886 33560 892
rect 29656 800 29684 886
rect 31588 800 31616 886
rect 33520 800 33548 886
rect 35452 800 35480 2382
rect 35728 2378 35756 5170
rect 35820 4282 35848 6174
rect 35992 6122 36044 6128
rect 35900 6112 35952 6118
rect 35900 6054 35952 6060
rect 35912 5778 35940 6054
rect 35900 5772 35952 5778
rect 35900 5714 35952 5720
rect 35808 4276 35860 4282
rect 35808 4218 35860 4224
rect 35912 4162 35940 5714
rect 36004 5234 36032 6122
rect 36084 5636 36136 5642
rect 36084 5578 36136 5584
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 35992 5024 36044 5030
rect 35992 4966 36044 4972
rect 36004 4282 36032 4966
rect 35992 4276 36044 4282
rect 35992 4218 36044 4224
rect 35820 4134 35940 4162
rect 35820 3602 35848 4134
rect 36096 3942 36124 5578
rect 36176 4820 36228 4826
rect 36176 4762 36228 4768
rect 36188 4622 36216 4762
rect 36176 4616 36228 4622
rect 36176 4558 36228 4564
rect 36266 4040 36322 4049
rect 36266 3975 36268 3984
rect 36320 3975 36322 3984
rect 36268 3946 36320 3952
rect 36084 3936 36136 3942
rect 36084 3878 36136 3884
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 35900 3392 35952 3398
rect 35900 3334 35952 3340
rect 35716 2372 35768 2378
rect 35716 2314 35768 2320
rect 35912 1873 35940 3334
rect 36372 2774 36400 12406
rect 36452 11008 36504 11014
rect 36452 10950 36504 10956
rect 36464 9994 36492 10950
rect 36556 10266 36584 23310
rect 37108 22710 37136 24006
rect 37096 22704 37148 22710
rect 37096 22646 37148 22652
rect 37568 21554 37596 25842
rect 37648 25696 37700 25702
rect 37648 25638 37700 25644
rect 37924 25696 37976 25702
rect 37924 25638 37976 25644
rect 37660 24682 37688 25638
rect 37648 24676 37700 24682
rect 37648 24618 37700 24624
rect 37556 21548 37608 21554
rect 37556 21490 37608 21496
rect 37186 19544 37242 19553
rect 37186 19479 37242 19488
rect 36820 18692 36872 18698
rect 36820 18634 36872 18640
rect 36832 18290 36860 18634
rect 37200 18426 37228 19479
rect 37464 19236 37516 19242
rect 37464 19178 37516 19184
rect 37476 18834 37504 19178
rect 37464 18828 37516 18834
rect 37464 18770 37516 18776
rect 37188 18420 37240 18426
rect 37188 18362 37240 18368
rect 36820 18284 36872 18290
rect 36820 18226 36872 18232
rect 37188 18284 37240 18290
rect 37188 18226 37240 18232
rect 36636 16584 36688 16590
rect 36636 16526 36688 16532
rect 36648 16114 36676 16526
rect 36636 16108 36688 16114
rect 36636 16050 36688 16056
rect 36728 15904 36780 15910
rect 36728 15846 36780 15852
rect 36740 15434 36768 15846
rect 36728 15428 36780 15434
rect 36728 15370 36780 15376
rect 36636 14816 36688 14822
rect 36636 14758 36688 14764
rect 36648 14385 36676 14758
rect 36634 14376 36690 14385
rect 36634 14311 36690 14320
rect 36636 14272 36688 14278
rect 36636 14214 36688 14220
rect 36728 14272 36780 14278
rect 36728 14214 36780 14220
rect 36648 14006 36676 14214
rect 36740 14074 36768 14214
rect 36728 14068 36780 14074
rect 36728 14010 36780 14016
rect 36636 14000 36688 14006
rect 36832 13954 36860 18226
rect 37200 17678 37228 18226
rect 37188 17672 37240 17678
rect 37188 17614 37240 17620
rect 37200 16114 37228 17614
rect 37372 17196 37424 17202
rect 37372 17138 37424 17144
rect 37188 16108 37240 16114
rect 37188 16050 37240 16056
rect 37096 15428 37148 15434
rect 37096 15370 37148 15376
rect 36636 13942 36688 13948
rect 36740 13926 36860 13954
rect 36636 10464 36688 10470
rect 36636 10406 36688 10412
rect 36544 10260 36596 10266
rect 36544 10202 36596 10208
rect 36452 9988 36504 9994
rect 36452 9930 36504 9936
rect 36544 9648 36596 9654
rect 36542 9616 36544 9625
rect 36596 9616 36598 9625
rect 36542 9551 36598 9560
rect 36544 6384 36596 6390
rect 36544 6326 36596 6332
rect 36556 4826 36584 6326
rect 36648 5370 36676 10406
rect 36740 8906 36768 13926
rect 36820 13864 36872 13870
rect 36820 13806 36872 13812
rect 36832 12434 36860 13806
rect 36832 12406 36952 12434
rect 36820 12096 36872 12102
rect 36820 12038 36872 12044
rect 36728 8900 36780 8906
rect 36728 8842 36780 8848
rect 36728 7200 36780 7206
rect 36728 7142 36780 7148
rect 36636 5364 36688 5370
rect 36636 5306 36688 5312
rect 36740 5030 36768 7142
rect 36832 6882 36860 12038
rect 36924 8945 36952 12406
rect 37108 11937 37136 15370
rect 37200 14414 37228 16050
rect 37280 15904 37332 15910
rect 37280 15846 37332 15852
rect 37188 14408 37240 14414
rect 37188 14350 37240 14356
rect 37292 13802 37320 15846
rect 37384 15570 37412 17138
rect 37556 16108 37608 16114
rect 37556 16050 37608 16056
rect 37372 15564 37424 15570
rect 37372 15506 37424 15512
rect 37372 14544 37424 14550
rect 37370 14512 37372 14521
rect 37424 14512 37426 14521
rect 37370 14447 37426 14456
rect 37280 13796 37332 13802
rect 37280 13738 37332 13744
rect 37372 13184 37424 13190
rect 37372 13126 37424 13132
rect 37186 12880 37242 12889
rect 37186 12815 37242 12824
rect 37200 12442 37228 12815
rect 37188 12436 37240 12442
rect 37384 12434 37412 13126
rect 37464 12844 37516 12850
rect 37464 12786 37516 12792
rect 37188 12378 37240 12384
rect 37292 12406 37412 12434
rect 37094 11928 37150 11937
rect 37094 11863 37150 11872
rect 37004 10192 37056 10198
rect 37004 10134 37056 10140
rect 36910 8936 36966 8945
rect 36910 8871 36966 8880
rect 36912 8424 36964 8430
rect 36912 8366 36964 8372
rect 36924 7546 36952 8366
rect 37016 7954 37044 10134
rect 37096 8900 37148 8906
rect 37096 8842 37148 8848
rect 37004 7948 37056 7954
rect 37004 7890 37056 7896
rect 36912 7540 36964 7546
rect 36912 7482 36964 7488
rect 36832 6854 37044 6882
rect 36820 6792 36872 6798
rect 36820 6734 36872 6740
rect 36910 6760 36966 6769
rect 36832 5778 36860 6734
rect 36910 6695 36966 6704
rect 36820 5772 36872 5778
rect 36820 5714 36872 5720
rect 36924 5370 36952 6695
rect 36912 5364 36964 5370
rect 36912 5306 36964 5312
rect 36818 5264 36874 5273
rect 36818 5199 36874 5208
rect 36728 5024 36780 5030
rect 36728 4966 36780 4972
rect 36544 4820 36596 4826
rect 36544 4762 36596 4768
rect 36636 3664 36688 3670
rect 36634 3632 36636 3641
rect 36688 3632 36690 3641
rect 36634 3567 36690 3576
rect 36832 3126 36860 5199
rect 36910 5128 36966 5137
rect 36910 5063 36912 5072
rect 36964 5063 36966 5072
rect 36912 5034 36964 5040
rect 37016 3602 37044 6854
rect 37108 6458 37136 8842
rect 37186 7712 37242 7721
rect 37186 7647 37242 7656
rect 37200 7546 37228 7647
rect 37188 7540 37240 7546
rect 37188 7482 37240 7488
rect 37096 6452 37148 6458
rect 37096 6394 37148 6400
rect 37292 5710 37320 12406
rect 37476 12306 37504 12786
rect 37464 12300 37516 12306
rect 37464 12242 37516 12248
rect 37464 11144 37516 11150
rect 37464 11086 37516 11092
rect 37372 10736 37424 10742
rect 37372 10678 37424 10684
rect 37384 8650 37412 10678
rect 37476 10062 37504 11086
rect 37568 10554 37596 16050
rect 37936 16046 37964 25638
rect 38948 25430 38976 28478
rect 39302 28354 39358 28478
rect 39394 27976 39450 27985
rect 39450 27934 39528 27962
rect 39394 27911 39450 27920
rect 39396 26376 39448 26382
rect 39396 26318 39448 26324
rect 39038 26140 39346 26149
rect 39038 26138 39044 26140
rect 39100 26138 39124 26140
rect 39180 26138 39204 26140
rect 39260 26138 39284 26140
rect 39340 26138 39346 26140
rect 39100 26086 39102 26138
rect 39282 26086 39284 26138
rect 39038 26084 39044 26086
rect 39100 26084 39124 26086
rect 39180 26084 39204 26086
rect 39260 26084 39284 26086
rect 39340 26084 39346 26086
rect 39038 26075 39346 26084
rect 39408 25945 39436 26318
rect 39500 25974 39528 27934
rect 39488 25968 39540 25974
rect 39394 25936 39450 25945
rect 39488 25910 39540 25916
rect 39394 25871 39450 25880
rect 38936 25424 38988 25430
rect 38936 25366 38988 25372
rect 39038 25052 39346 25061
rect 39038 25050 39044 25052
rect 39100 25050 39124 25052
rect 39180 25050 39204 25052
rect 39260 25050 39284 25052
rect 39340 25050 39346 25052
rect 39100 24998 39102 25050
rect 39282 24998 39284 25050
rect 39038 24996 39044 24998
rect 39100 24996 39124 24998
rect 39180 24996 39204 24998
rect 39260 24996 39284 24998
rect 39340 24996 39346 24998
rect 39038 24987 39346 24996
rect 39396 24812 39448 24818
rect 39396 24754 39448 24760
rect 38292 24744 38344 24750
rect 38292 24686 38344 24692
rect 38304 23798 38332 24686
rect 39408 24585 39436 24754
rect 39394 24576 39450 24585
rect 39394 24511 39450 24520
rect 39038 23964 39346 23973
rect 39038 23962 39044 23964
rect 39100 23962 39124 23964
rect 39180 23962 39204 23964
rect 39260 23962 39284 23964
rect 39340 23962 39346 23964
rect 39100 23910 39102 23962
rect 39282 23910 39284 23962
rect 39038 23908 39044 23910
rect 39100 23908 39124 23910
rect 39180 23908 39204 23910
rect 39260 23908 39284 23910
rect 39340 23908 39346 23910
rect 39038 23899 39346 23908
rect 38292 23792 38344 23798
rect 38292 23734 38344 23740
rect 39038 22876 39346 22885
rect 39038 22874 39044 22876
rect 39100 22874 39124 22876
rect 39180 22874 39204 22876
rect 39260 22874 39284 22876
rect 39340 22874 39346 22876
rect 39100 22822 39102 22874
rect 39282 22822 39284 22874
rect 39038 22820 39044 22822
rect 39100 22820 39124 22822
rect 39180 22820 39204 22822
rect 39260 22820 39284 22822
rect 39340 22820 39346 22822
rect 39038 22811 39346 22820
rect 39038 21788 39346 21797
rect 39038 21786 39044 21788
rect 39100 21786 39124 21788
rect 39180 21786 39204 21788
rect 39260 21786 39284 21788
rect 39340 21786 39346 21788
rect 39100 21734 39102 21786
rect 39282 21734 39284 21786
rect 39038 21732 39044 21734
rect 39100 21732 39124 21734
rect 39180 21732 39204 21734
rect 39260 21732 39284 21734
rect 39340 21732 39346 21734
rect 39038 21723 39346 21732
rect 38476 20868 38528 20874
rect 38476 20810 38528 20816
rect 39396 20868 39448 20874
rect 39396 20810 39448 20816
rect 38488 19961 38516 20810
rect 39038 20700 39346 20709
rect 39038 20698 39044 20700
rect 39100 20698 39124 20700
rect 39180 20698 39204 20700
rect 39260 20698 39284 20700
rect 39340 20698 39346 20700
rect 39100 20646 39102 20698
rect 39282 20646 39284 20698
rect 39038 20644 39044 20646
rect 39100 20644 39124 20646
rect 39180 20644 39204 20646
rect 39260 20644 39284 20646
rect 39340 20644 39346 20646
rect 39038 20635 39346 20644
rect 39408 20505 39436 20810
rect 39394 20496 39450 20505
rect 39394 20431 39450 20440
rect 38474 19952 38530 19961
rect 38474 19887 38530 19896
rect 39038 19612 39346 19621
rect 39038 19610 39044 19612
rect 39100 19610 39124 19612
rect 39180 19610 39204 19612
rect 39260 19610 39284 19612
rect 39340 19610 39346 19612
rect 39100 19558 39102 19610
rect 39282 19558 39284 19610
rect 39038 19556 39044 19558
rect 39100 19556 39124 19558
rect 39180 19556 39204 19558
rect 39260 19556 39284 19558
rect 39340 19556 39346 19558
rect 39038 19547 39346 19556
rect 39038 18524 39346 18533
rect 39038 18522 39044 18524
rect 39100 18522 39124 18524
rect 39180 18522 39204 18524
rect 39260 18522 39284 18524
rect 39340 18522 39346 18524
rect 39100 18470 39102 18522
rect 39282 18470 39284 18522
rect 39038 18468 39044 18470
rect 39100 18468 39124 18470
rect 39180 18468 39204 18470
rect 39260 18468 39284 18470
rect 39340 18468 39346 18470
rect 39038 18459 39346 18468
rect 39038 17436 39346 17445
rect 39038 17434 39044 17436
rect 39100 17434 39124 17436
rect 39180 17434 39204 17436
rect 39260 17434 39284 17436
rect 39340 17434 39346 17436
rect 39100 17382 39102 17434
rect 39282 17382 39284 17434
rect 39038 17380 39044 17382
rect 39100 17380 39124 17382
rect 39180 17380 39204 17382
rect 39260 17380 39284 17382
rect 39340 17380 39346 17382
rect 39038 17371 39346 17380
rect 38568 17332 38620 17338
rect 38568 17274 38620 17280
rect 38476 16176 38528 16182
rect 38476 16118 38528 16124
rect 37924 16040 37976 16046
rect 37924 15982 37976 15988
rect 37936 15502 37964 15982
rect 37924 15496 37976 15502
rect 37924 15438 37976 15444
rect 38488 15094 38516 16118
rect 38476 15088 38528 15094
rect 38476 15030 38528 15036
rect 37832 15020 37884 15026
rect 37832 14962 37884 14968
rect 37844 13870 37872 14962
rect 38108 14408 38160 14414
rect 38108 14350 38160 14356
rect 38120 13938 38148 14350
rect 38108 13932 38160 13938
rect 38108 13874 38160 13880
rect 37832 13864 37884 13870
rect 37832 13806 37884 13812
rect 37740 13184 37792 13190
rect 37740 13126 37792 13132
rect 37648 11076 37700 11082
rect 37648 11018 37700 11024
rect 37660 10713 37688 11018
rect 37752 11014 37780 13126
rect 37844 12850 37872 13806
rect 37832 12844 37884 12850
rect 37832 12786 37884 12792
rect 37740 11008 37792 11014
rect 37740 10950 37792 10956
rect 37646 10704 37702 10713
rect 37844 10674 37872 12786
rect 38016 12232 38068 12238
rect 38016 12174 38068 12180
rect 38028 11762 38056 12174
rect 38016 11756 38068 11762
rect 38016 11698 38068 11704
rect 38120 11150 38148 13874
rect 38200 13728 38252 13734
rect 38200 13670 38252 13676
rect 38212 13258 38240 13670
rect 38384 13320 38436 13326
rect 38384 13262 38436 13268
rect 38200 13252 38252 13258
rect 38200 13194 38252 13200
rect 38292 12640 38344 12646
rect 38292 12582 38344 12588
rect 38108 11144 38160 11150
rect 38108 11086 38160 11092
rect 37646 10639 37702 10648
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 38016 10668 38068 10674
rect 38068 10628 38148 10656
rect 38016 10610 38068 10616
rect 37568 10526 37780 10554
rect 37648 10464 37700 10470
rect 37648 10406 37700 10412
rect 37464 10056 37516 10062
rect 37464 9998 37516 10004
rect 37476 9586 37504 9998
rect 37556 9920 37608 9926
rect 37556 9862 37608 9868
rect 37464 9580 37516 9586
rect 37464 9522 37516 9528
rect 37568 8906 37596 9862
rect 37556 8900 37608 8906
rect 37556 8842 37608 8848
rect 37384 8622 37504 8650
rect 37370 8528 37426 8537
rect 37370 8463 37426 8472
rect 37384 7886 37412 8463
rect 37372 7880 37424 7886
rect 37372 7822 37424 7828
rect 37372 6724 37424 6730
rect 37372 6666 37424 6672
rect 37280 5704 37332 5710
rect 37280 5646 37332 5652
rect 37188 5568 37240 5574
rect 37188 5510 37240 5516
rect 37200 4826 37228 5510
rect 37188 4820 37240 4826
rect 37188 4762 37240 4768
rect 37188 4616 37240 4622
rect 37240 4564 37320 4570
rect 37188 4558 37320 4564
rect 37096 4548 37148 4554
rect 37200 4542 37320 4558
rect 37096 4490 37148 4496
rect 37004 3596 37056 3602
rect 37004 3538 37056 3544
rect 37108 3534 37136 4490
rect 37292 4146 37320 4542
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 37292 3738 37320 4082
rect 37280 3732 37332 3738
rect 37280 3674 37332 3680
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 36820 3120 36872 3126
rect 36820 3062 36872 3068
rect 37108 3058 37136 3470
rect 37280 3392 37332 3398
rect 37280 3334 37332 3340
rect 37096 3052 37148 3058
rect 37096 2994 37148 3000
rect 36820 2984 36872 2990
rect 36818 2952 36820 2961
rect 36872 2952 36874 2961
rect 36818 2887 36874 2896
rect 36004 2746 36400 2774
rect 36004 2106 36032 2746
rect 36636 2304 36688 2310
rect 36636 2246 36688 2252
rect 35992 2100 36044 2106
rect 35992 2042 36044 2048
rect 35898 1864 35954 1873
rect 35898 1799 35954 1808
rect 36648 950 36676 2246
rect 37292 2009 37320 3334
rect 37278 2000 37334 2009
rect 37278 1935 37334 1944
rect 37384 1358 37412 6666
rect 37476 5370 37504 8622
rect 37554 8120 37610 8129
rect 37554 8055 37610 8064
rect 37464 5364 37516 5370
rect 37464 5306 37516 5312
rect 37464 5228 37516 5234
rect 37464 5170 37516 5176
rect 37476 4554 37504 5170
rect 37568 4622 37596 8055
rect 37556 4616 37608 4622
rect 37556 4558 37608 4564
rect 37464 4548 37516 4554
rect 37464 4490 37516 4496
rect 37476 3194 37504 4490
rect 37660 4185 37688 10406
rect 37752 8129 37780 10526
rect 38120 9586 38148 10628
rect 38200 10464 38252 10470
rect 38200 10406 38252 10412
rect 38212 10169 38240 10406
rect 38198 10160 38254 10169
rect 38198 10095 38254 10104
rect 38108 9580 38160 9586
rect 38108 9522 38160 9528
rect 37924 9512 37976 9518
rect 37924 9454 37976 9460
rect 37936 8634 37964 9454
rect 37924 8628 37976 8634
rect 37924 8570 37976 8576
rect 37832 8492 37884 8498
rect 37832 8434 37884 8440
rect 37738 8120 37794 8129
rect 37738 8055 37794 8064
rect 37740 8016 37792 8022
rect 37738 7984 37740 7993
rect 37792 7984 37794 7993
rect 37738 7919 37794 7928
rect 37740 7336 37792 7342
rect 37740 7278 37792 7284
rect 37752 6866 37780 7278
rect 37740 6860 37792 6866
rect 37740 6802 37792 6808
rect 37844 6662 37872 8434
rect 37832 6656 37884 6662
rect 37832 6598 37884 6604
rect 37936 6338 37964 8570
rect 37844 6310 37964 6338
rect 37844 5302 37872 6310
rect 37924 6248 37976 6254
rect 37924 6190 37976 6196
rect 37936 5930 37964 6190
rect 37936 5914 38056 5930
rect 37936 5908 38068 5914
rect 37936 5902 38016 5908
rect 38016 5850 38068 5856
rect 37832 5296 37884 5302
rect 37832 5238 37884 5244
rect 38120 5234 38148 9522
rect 38200 9376 38252 9382
rect 38200 9318 38252 9324
rect 38212 8401 38240 9318
rect 38198 8392 38254 8401
rect 38198 8327 38254 8336
rect 38108 5228 38160 5234
rect 38108 5170 38160 5176
rect 37646 4176 37702 4185
rect 38120 4146 38148 5170
rect 38304 4486 38332 12582
rect 38396 12238 38424 13262
rect 38384 12232 38436 12238
rect 38384 12174 38436 12180
rect 38396 10674 38424 12174
rect 38384 10668 38436 10674
rect 38384 10610 38436 10616
rect 38396 5710 38424 10610
rect 38580 9178 38608 17274
rect 38658 17096 38714 17105
rect 38658 17031 38660 17040
rect 38712 17031 38714 17040
rect 38660 17002 38712 17008
rect 39038 16348 39346 16357
rect 39038 16346 39044 16348
rect 39100 16346 39124 16348
rect 39180 16346 39204 16348
rect 39260 16346 39284 16348
rect 39340 16346 39346 16348
rect 39100 16294 39102 16346
rect 39282 16294 39284 16346
rect 39038 16292 39044 16294
rect 39100 16292 39124 16294
rect 39180 16292 39204 16294
rect 39260 16292 39284 16294
rect 39340 16292 39346 16294
rect 39038 16283 39346 16292
rect 39038 15260 39346 15269
rect 39038 15258 39044 15260
rect 39100 15258 39124 15260
rect 39180 15258 39204 15260
rect 39260 15258 39284 15260
rect 39340 15258 39346 15260
rect 39100 15206 39102 15258
rect 39282 15206 39284 15258
rect 39038 15204 39044 15206
rect 39100 15204 39124 15206
rect 39180 15204 39204 15206
rect 39260 15204 39284 15206
rect 39340 15204 39346 15206
rect 39038 15195 39346 15204
rect 38658 15056 38714 15065
rect 38658 14991 38660 15000
rect 38712 14991 38714 15000
rect 38660 14962 38712 14968
rect 39038 14172 39346 14181
rect 39038 14170 39044 14172
rect 39100 14170 39124 14172
rect 39180 14170 39204 14172
rect 39260 14170 39284 14172
rect 39340 14170 39346 14172
rect 39100 14118 39102 14170
rect 39282 14118 39284 14170
rect 39038 14116 39044 14118
rect 39100 14116 39124 14118
rect 39180 14116 39204 14118
rect 39260 14116 39284 14118
rect 39340 14116 39346 14118
rect 39038 14107 39346 14116
rect 39396 13252 39448 13258
rect 39396 13194 39448 13200
rect 39038 13084 39346 13093
rect 39038 13082 39044 13084
rect 39100 13082 39124 13084
rect 39180 13082 39204 13084
rect 39260 13082 39284 13084
rect 39340 13082 39346 13084
rect 39100 13030 39102 13082
rect 39282 13030 39284 13082
rect 39038 13028 39044 13030
rect 39100 13028 39124 13030
rect 39180 13028 39204 13030
rect 39260 13028 39284 13030
rect 39340 13028 39346 13030
rect 39038 13019 39346 13028
rect 39408 12889 39436 13194
rect 39394 12880 39450 12889
rect 39394 12815 39450 12824
rect 39038 11996 39346 12005
rect 39038 11994 39044 11996
rect 39100 11994 39124 11996
rect 39180 11994 39204 11996
rect 39260 11994 39284 11996
rect 39340 11994 39346 11996
rect 39100 11942 39102 11994
rect 39282 11942 39284 11994
rect 39038 11940 39044 11942
rect 39100 11940 39124 11942
rect 39180 11940 39204 11942
rect 39260 11940 39284 11942
rect 39340 11940 39346 11942
rect 39038 11931 39346 11940
rect 39394 11112 39450 11121
rect 39394 11047 39396 11056
rect 39448 11047 39450 11056
rect 39396 11018 39448 11024
rect 39038 10908 39346 10917
rect 39038 10906 39044 10908
rect 39100 10906 39124 10908
rect 39180 10906 39204 10908
rect 39260 10906 39284 10908
rect 39340 10906 39346 10908
rect 39100 10854 39102 10906
rect 39282 10854 39284 10906
rect 39038 10852 39044 10854
rect 39100 10852 39124 10854
rect 39180 10852 39204 10854
rect 39260 10852 39284 10854
rect 39340 10852 39346 10854
rect 39038 10843 39346 10852
rect 39396 10056 39448 10062
rect 39396 9998 39448 10004
rect 39038 9820 39346 9829
rect 39038 9818 39044 9820
rect 39100 9818 39124 9820
rect 39180 9818 39204 9820
rect 39260 9818 39284 9820
rect 39340 9818 39346 9820
rect 39100 9766 39102 9818
rect 39282 9766 39284 9818
rect 39038 9764 39044 9766
rect 39100 9764 39124 9766
rect 39180 9764 39204 9766
rect 39260 9764 39284 9766
rect 39340 9764 39346 9766
rect 39038 9755 39346 9764
rect 39408 9625 39436 9998
rect 39394 9616 39450 9625
rect 39394 9551 39450 9560
rect 38568 9172 38620 9178
rect 38568 9114 38620 9120
rect 38580 6746 38608 9114
rect 39038 8732 39346 8741
rect 39038 8730 39044 8732
rect 39100 8730 39124 8732
rect 39180 8730 39204 8732
rect 39260 8730 39284 8732
rect 39340 8730 39346 8732
rect 39100 8678 39102 8730
rect 39282 8678 39284 8730
rect 39038 8676 39044 8678
rect 39100 8676 39124 8678
rect 39180 8676 39204 8678
rect 39260 8676 39284 8678
rect 39340 8676 39346 8678
rect 39038 8667 39346 8676
rect 38660 7812 38712 7818
rect 38660 7754 38712 7760
rect 38672 7449 38700 7754
rect 39038 7644 39346 7653
rect 39038 7642 39044 7644
rect 39100 7642 39124 7644
rect 39180 7642 39204 7644
rect 39260 7642 39284 7644
rect 39340 7642 39346 7644
rect 39100 7590 39102 7642
rect 39282 7590 39284 7642
rect 39038 7588 39044 7590
rect 39100 7588 39124 7590
rect 39180 7588 39204 7590
rect 39260 7588 39284 7590
rect 39340 7588 39346 7590
rect 39038 7579 39346 7588
rect 38658 7440 38714 7449
rect 38658 7375 38714 7384
rect 38488 6718 38608 6746
rect 38488 6458 38516 6718
rect 38568 6656 38620 6662
rect 38568 6598 38620 6604
rect 38476 6452 38528 6458
rect 38476 6394 38528 6400
rect 38384 5704 38436 5710
rect 38384 5646 38436 5652
rect 38396 4554 38424 5646
rect 38384 4548 38436 4554
rect 38384 4490 38436 4496
rect 38292 4480 38344 4486
rect 38292 4422 38344 4428
rect 37646 4111 37702 4120
rect 38108 4140 38160 4146
rect 38108 4082 38160 4088
rect 38200 3936 38252 3942
rect 38200 3878 38252 3884
rect 37464 3188 37516 3194
rect 37464 3130 37516 3136
rect 37556 2848 37608 2854
rect 37556 2790 37608 2796
rect 37568 1970 37596 2790
rect 37648 2304 37700 2310
rect 37648 2246 37700 2252
rect 37556 1964 37608 1970
rect 37556 1906 37608 1912
rect 37372 1352 37424 1358
rect 37372 1294 37424 1300
rect 37660 950 37688 2246
rect 38212 1737 38240 3878
rect 38474 2408 38530 2417
rect 38474 2343 38476 2352
rect 38528 2343 38530 2352
rect 38476 2314 38528 2320
rect 38198 1728 38254 1737
rect 38198 1663 38254 1672
rect 38580 1290 38608 6598
rect 39038 6556 39346 6565
rect 39038 6554 39044 6556
rect 39100 6554 39124 6556
rect 39180 6554 39204 6556
rect 39260 6554 39284 6556
rect 39340 6554 39346 6556
rect 39100 6502 39102 6554
rect 39282 6502 39284 6554
rect 39038 6500 39044 6502
rect 39100 6500 39124 6502
rect 39180 6500 39204 6502
rect 39260 6500 39284 6502
rect 39340 6500 39346 6502
rect 39038 6491 39346 6500
rect 39038 5468 39346 5477
rect 39038 5466 39044 5468
rect 39100 5466 39124 5468
rect 39180 5466 39204 5468
rect 39260 5466 39284 5468
rect 39340 5466 39346 5468
rect 39100 5414 39102 5466
rect 39282 5414 39284 5466
rect 39038 5412 39044 5414
rect 39100 5412 39124 5414
rect 39180 5412 39204 5414
rect 39260 5412 39284 5414
rect 39340 5412 39346 5414
rect 39038 5403 39346 5412
rect 39038 4380 39346 4389
rect 39038 4378 39044 4380
rect 39100 4378 39124 4380
rect 39180 4378 39204 4380
rect 39260 4378 39284 4380
rect 39340 4378 39346 4380
rect 39100 4326 39102 4378
rect 39282 4326 39284 4378
rect 39038 4324 39044 4326
rect 39100 4324 39124 4326
rect 39180 4324 39204 4326
rect 39260 4324 39284 4326
rect 39340 4324 39346 4326
rect 39038 4315 39346 4324
rect 38658 3496 38714 3505
rect 38658 3431 38660 3440
rect 38712 3431 38714 3440
rect 38660 3402 38712 3408
rect 39038 3292 39346 3301
rect 39038 3290 39044 3292
rect 39100 3290 39124 3292
rect 39180 3290 39204 3292
rect 39260 3290 39284 3292
rect 39340 3290 39346 3292
rect 39100 3238 39102 3290
rect 39282 3238 39284 3290
rect 39038 3236 39044 3238
rect 39100 3236 39124 3238
rect 39180 3236 39204 3238
rect 39260 3236 39284 3238
rect 39340 3236 39346 3238
rect 39038 3227 39346 3236
rect 39396 2916 39448 2922
rect 39396 2858 39448 2864
rect 38660 2372 38712 2378
rect 38660 2314 38712 2320
rect 38672 2009 38700 2314
rect 39038 2204 39346 2213
rect 39038 2202 39044 2204
rect 39100 2202 39124 2204
rect 39180 2202 39204 2204
rect 39260 2202 39284 2204
rect 39340 2202 39346 2204
rect 39100 2150 39102 2202
rect 39282 2150 39284 2202
rect 39038 2148 39044 2150
rect 39100 2148 39124 2150
rect 39180 2148 39204 2150
rect 39260 2148 39284 2150
rect 39340 2148 39346 2150
rect 39038 2139 39346 2148
rect 38658 2000 38714 2009
rect 38658 1935 38714 1944
rect 38568 1284 38620 1290
rect 38568 1226 38620 1232
rect 36636 944 36688 950
rect 36636 886 36688 892
rect 36728 944 36780 950
rect 36728 886 36780 892
rect 37648 944 37700 950
rect 37648 886 37700 892
rect 36740 800 36768 886
rect 13924 734 14136 762
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 17406 0 17462 800
rect 19338 0 19394 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 31574 0 31630 800
rect 33506 0 33562 800
rect 35438 0 35494 800
rect 36726 0 36782 800
rect 38658 0 38714 800
rect 39408 105 39436 2858
rect 39394 96 39450 105
rect 39394 31 39450 40
<< via2 >>
rect 1030 27920 1086 27976
rect 938 25880 994 25936
rect 5717 26682 5773 26684
rect 5797 26682 5853 26684
rect 5877 26682 5933 26684
rect 5957 26682 6013 26684
rect 5717 26630 5763 26682
rect 5763 26630 5773 26682
rect 5797 26630 5827 26682
rect 5827 26630 5839 26682
rect 5839 26630 5853 26682
rect 5877 26630 5891 26682
rect 5891 26630 5903 26682
rect 5903 26630 5933 26682
rect 5957 26630 5967 26682
rect 5967 26630 6013 26682
rect 5717 26628 5773 26630
rect 5797 26628 5853 26630
rect 5877 26628 5933 26630
rect 5957 26628 6013 26630
rect 3054 26308 3110 26344
rect 3054 26288 3056 26308
rect 3056 26288 3108 26308
rect 3108 26288 3110 26308
rect 7930 26308 7986 26344
rect 7930 26288 7932 26308
rect 7932 26288 7984 26308
rect 7984 26288 7986 26308
rect 938 23840 994 23896
rect 938 22480 994 22536
rect 938 20440 994 20496
rect 938 18400 994 18456
rect 938 16360 994 16416
rect 938 15000 994 15056
rect 1674 13776 1730 13832
rect 938 12960 994 13016
rect 2042 15544 2098 15600
rect 5717 25594 5773 25596
rect 5797 25594 5853 25596
rect 5877 25594 5933 25596
rect 5957 25594 6013 25596
rect 5717 25542 5763 25594
rect 5763 25542 5773 25594
rect 5797 25542 5827 25594
rect 5827 25542 5839 25594
rect 5839 25542 5853 25594
rect 5877 25542 5891 25594
rect 5891 25542 5903 25594
rect 5903 25542 5933 25594
rect 5957 25542 5967 25594
rect 5967 25542 6013 25594
rect 5717 25540 5773 25542
rect 5797 25540 5853 25542
rect 5877 25540 5933 25542
rect 5957 25540 6013 25542
rect 5717 24506 5773 24508
rect 5797 24506 5853 24508
rect 5877 24506 5933 24508
rect 5957 24506 6013 24508
rect 5717 24454 5763 24506
rect 5763 24454 5773 24506
rect 5797 24454 5827 24506
rect 5827 24454 5839 24506
rect 5839 24454 5853 24506
rect 5877 24454 5891 24506
rect 5891 24454 5903 24506
rect 5903 24454 5933 24506
rect 5957 24454 5967 24506
rect 5967 24454 6013 24506
rect 5717 24452 5773 24454
rect 5797 24452 5853 24454
rect 5877 24452 5933 24454
rect 5957 24452 6013 24454
rect 1858 11192 1914 11248
rect 938 10920 994 10976
rect 938 8880 994 8936
rect 938 7520 994 7576
rect 1030 5480 1086 5536
rect 938 3440 994 3496
rect 1766 9424 1822 9480
rect 2778 16632 2834 16688
rect 2686 15136 2742 15192
rect 2226 9988 2282 10024
rect 2226 9968 2228 9988
rect 2228 9968 2280 9988
rect 2280 9968 2282 9988
rect 1858 3596 1914 3632
rect 1858 3576 1860 3596
rect 1860 3576 1912 3596
rect 1912 3576 1914 3596
rect 1858 3168 1914 3224
rect 2778 12144 2834 12200
rect 2594 9696 2650 9752
rect 2778 7928 2834 7984
rect 2778 7112 2834 7168
rect 2686 5616 2742 5672
rect 3054 15308 3056 15328
rect 3056 15308 3108 15328
rect 3108 15308 3110 15328
rect 3054 15272 3110 15308
rect 3422 17584 3478 17640
rect 3330 13268 3332 13288
rect 3332 13268 3384 13288
rect 3384 13268 3386 13288
rect 3330 13232 3386 13268
rect 2778 4256 2834 4312
rect 3054 6840 3110 6896
rect 3146 6432 3202 6488
rect 3514 12144 3570 12200
rect 3422 8472 3478 8528
rect 4342 15408 4398 15464
rect 4526 15816 4582 15872
rect 5717 23418 5773 23420
rect 5797 23418 5853 23420
rect 5877 23418 5933 23420
rect 5957 23418 6013 23420
rect 5717 23366 5763 23418
rect 5763 23366 5773 23418
rect 5797 23366 5827 23418
rect 5827 23366 5839 23418
rect 5839 23366 5853 23418
rect 5877 23366 5891 23418
rect 5891 23366 5903 23418
rect 5903 23366 5933 23418
rect 5957 23366 5967 23418
rect 5967 23366 6013 23418
rect 5717 23364 5773 23366
rect 5797 23364 5853 23366
rect 5877 23364 5933 23366
rect 5957 23364 6013 23366
rect 5717 22330 5773 22332
rect 5797 22330 5853 22332
rect 5877 22330 5933 22332
rect 5957 22330 6013 22332
rect 5717 22278 5763 22330
rect 5763 22278 5773 22330
rect 5797 22278 5827 22330
rect 5827 22278 5839 22330
rect 5839 22278 5853 22330
rect 5877 22278 5891 22330
rect 5891 22278 5903 22330
rect 5903 22278 5933 22330
rect 5957 22278 5967 22330
rect 5967 22278 6013 22330
rect 5717 22276 5773 22278
rect 5797 22276 5853 22278
rect 5877 22276 5933 22278
rect 5957 22276 6013 22278
rect 5717 21242 5773 21244
rect 5797 21242 5853 21244
rect 5877 21242 5933 21244
rect 5957 21242 6013 21244
rect 5717 21190 5763 21242
rect 5763 21190 5773 21242
rect 5797 21190 5827 21242
rect 5827 21190 5839 21242
rect 5839 21190 5853 21242
rect 5877 21190 5891 21242
rect 5891 21190 5903 21242
rect 5903 21190 5933 21242
rect 5957 21190 5967 21242
rect 5967 21190 6013 21242
rect 5717 21188 5773 21190
rect 5797 21188 5853 21190
rect 5877 21188 5933 21190
rect 5957 21188 6013 21190
rect 5717 20154 5773 20156
rect 5797 20154 5853 20156
rect 5877 20154 5933 20156
rect 5957 20154 6013 20156
rect 5717 20102 5763 20154
rect 5763 20102 5773 20154
rect 5797 20102 5827 20154
rect 5827 20102 5839 20154
rect 5839 20102 5853 20154
rect 5877 20102 5891 20154
rect 5891 20102 5903 20154
rect 5903 20102 5933 20154
rect 5957 20102 5967 20154
rect 5967 20102 6013 20154
rect 5717 20100 5773 20102
rect 5797 20100 5853 20102
rect 5877 20100 5933 20102
rect 5957 20100 6013 20102
rect 5717 19066 5773 19068
rect 5797 19066 5853 19068
rect 5877 19066 5933 19068
rect 5957 19066 6013 19068
rect 5717 19014 5763 19066
rect 5763 19014 5773 19066
rect 5797 19014 5827 19066
rect 5827 19014 5839 19066
rect 5839 19014 5853 19066
rect 5877 19014 5891 19066
rect 5891 19014 5903 19066
rect 5903 19014 5933 19066
rect 5957 19014 5967 19066
rect 5967 19014 6013 19066
rect 5717 19012 5773 19014
rect 5797 19012 5853 19014
rect 5877 19012 5933 19014
rect 5957 19012 6013 19014
rect 5170 17040 5226 17096
rect 4802 15272 4858 15328
rect 4894 15000 4950 15056
rect 4986 14456 5042 14512
rect 3606 7656 3662 7712
rect 3514 6432 3570 6488
rect 3698 5616 3754 5672
rect 3514 3596 3570 3632
rect 3514 3576 3516 3596
rect 3516 3576 3568 3596
rect 3568 3576 3570 3596
rect 4066 8608 4122 8664
rect 4066 7520 4122 7576
rect 4894 11600 4950 11656
rect 4342 7248 4398 7304
rect 4618 8608 4674 8664
rect 4526 6840 4582 6896
rect 3974 3984 4030 4040
rect 1398 1400 1454 1456
rect 4342 5752 4398 5808
rect 4526 5480 4582 5536
rect 4526 4120 4582 4176
rect 4802 7404 4858 7440
rect 4802 7384 4804 7404
rect 4804 7384 4856 7404
rect 4856 7384 4858 7404
rect 5354 17040 5410 17096
rect 5717 17978 5773 17980
rect 5797 17978 5853 17980
rect 5877 17978 5933 17980
rect 5957 17978 6013 17980
rect 5717 17926 5763 17978
rect 5763 17926 5773 17978
rect 5797 17926 5827 17978
rect 5827 17926 5839 17978
rect 5839 17926 5853 17978
rect 5877 17926 5891 17978
rect 5891 17926 5903 17978
rect 5903 17926 5933 17978
rect 5957 17926 5967 17978
rect 5967 17926 6013 17978
rect 5717 17924 5773 17926
rect 5797 17924 5853 17926
rect 5877 17924 5933 17926
rect 5957 17924 6013 17926
rect 5717 16890 5773 16892
rect 5797 16890 5853 16892
rect 5877 16890 5933 16892
rect 5957 16890 6013 16892
rect 5717 16838 5763 16890
rect 5763 16838 5773 16890
rect 5797 16838 5827 16890
rect 5827 16838 5839 16890
rect 5839 16838 5853 16890
rect 5877 16838 5891 16890
rect 5891 16838 5903 16890
rect 5903 16838 5933 16890
rect 5957 16838 5967 16890
rect 5967 16838 6013 16890
rect 5717 16836 5773 16838
rect 5797 16836 5853 16838
rect 5877 16836 5933 16838
rect 5957 16836 6013 16838
rect 5717 15802 5773 15804
rect 5797 15802 5853 15804
rect 5877 15802 5933 15804
rect 5957 15802 6013 15804
rect 5717 15750 5763 15802
rect 5763 15750 5773 15802
rect 5797 15750 5827 15802
rect 5827 15750 5839 15802
rect 5839 15750 5853 15802
rect 5877 15750 5891 15802
rect 5891 15750 5903 15802
rect 5903 15750 5933 15802
rect 5957 15750 5967 15802
rect 5967 15750 6013 15802
rect 5717 15748 5773 15750
rect 5797 15748 5853 15750
rect 5877 15748 5933 15750
rect 5957 15748 6013 15750
rect 5717 14714 5773 14716
rect 5797 14714 5853 14716
rect 5877 14714 5933 14716
rect 5957 14714 6013 14716
rect 5717 14662 5763 14714
rect 5763 14662 5773 14714
rect 5797 14662 5827 14714
rect 5827 14662 5839 14714
rect 5839 14662 5853 14714
rect 5877 14662 5891 14714
rect 5891 14662 5903 14714
rect 5903 14662 5933 14714
rect 5957 14662 5967 14714
rect 5967 14662 6013 14714
rect 5717 14660 5773 14662
rect 5797 14660 5853 14662
rect 5877 14660 5933 14662
rect 5957 14660 6013 14662
rect 5717 13626 5773 13628
rect 5797 13626 5853 13628
rect 5877 13626 5933 13628
rect 5957 13626 6013 13628
rect 5717 13574 5763 13626
rect 5763 13574 5773 13626
rect 5797 13574 5827 13626
rect 5827 13574 5839 13626
rect 5839 13574 5853 13626
rect 5877 13574 5891 13626
rect 5891 13574 5903 13626
rect 5903 13574 5933 13626
rect 5957 13574 5967 13626
rect 5967 13574 6013 13626
rect 5717 13572 5773 13574
rect 5797 13572 5853 13574
rect 5877 13572 5933 13574
rect 5957 13572 6013 13574
rect 5262 12588 5264 12608
rect 5264 12588 5316 12608
rect 5316 12588 5318 12608
rect 5262 12552 5318 12588
rect 6918 18264 6974 18320
rect 6642 15272 6698 15328
rect 5717 12538 5773 12540
rect 5797 12538 5853 12540
rect 5877 12538 5933 12540
rect 5957 12538 6013 12540
rect 5717 12486 5763 12538
rect 5763 12486 5773 12538
rect 5797 12486 5827 12538
rect 5827 12486 5839 12538
rect 5839 12486 5853 12538
rect 5877 12486 5891 12538
rect 5891 12486 5903 12538
rect 5903 12486 5933 12538
rect 5957 12486 5967 12538
rect 5967 12486 6013 12538
rect 5717 12484 5773 12486
rect 5797 12484 5853 12486
rect 5877 12484 5933 12486
rect 5957 12484 6013 12486
rect 7102 14456 7158 14512
rect 6734 13912 6790 13968
rect 6642 13676 6644 13696
rect 6644 13676 6696 13696
rect 6696 13676 6698 13696
rect 6642 13640 6698 13676
rect 5078 11600 5134 11656
rect 4894 7248 4950 7304
rect 5446 10512 5502 10568
rect 5814 11636 5816 11656
rect 5816 11636 5868 11656
rect 5868 11636 5870 11656
rect 5814 11600 5870 11636
rect 5717 11450 5773 11452
rect 5797 11450 5853 11452
rect 5877 11450 5933 11452
rect 5957 11450 6013 11452
rect 5717 11398 5763 11450
rect 5763 11398 5773 11450
rect 5797 11398 5827 11450
rect 5827 11398 5839 11450
rect 5839 11398 5853 11450
rect 5877 11398 5891 11450
rect 5891 11398 5903 11450
rect 5903 11398 5933 11450
rect 5957 11398 5967 11450
rect 5967 11398 6013 11450
rect 5717 11396 5773 11398
rect 5797 11396 5853 11398
rect 5877 11396 5933 11398
rect 5957 11396 6013 11398
rect 5722 10684 5724 10704
rect 5724 10684 5776 10704
rect 5776 10684 5778 10704
rect 5722 10648 5778 10684
rect 5717 10362 5773 10364
rect 5797 10362 5853 10364
rect 5877 10362 5933 10364
rect 5957 10362 6013 10364
rect 5717 10310 5763 10362
rect 5763 10310 5773 10362
rect 5797 10310 5827 10362
rect 5827 10310 5839 10362
rect 5839 10310 5853 10362
rect 5877 10310 5891 10362
rect 5891 10310 5903 10362
rect 5903 10310 5933 10362
rect 5957 10310 5967 10362
rect 5967 10310 6013 10362
rect 5717 10308 5773 10310
rect 5797 10308 5853 10310
rect 5877 10308 5933 10310
rect 5957 10308 6013 10310
rect 5446 8472 5502 8528
rect 5170 6296 5226 6352
rect 5354 6568 5410 6624
rect 5717 9274 5773 9276
rect 5797 9274 5853 9276
rect 5877 9274 5933 9276
rect 5957 9274 6013 9276
rect 5717 9222 5763 9274
rect 5763 9222 5773 9274
rect 5797 9222 5827 9274
rect 5827 9222 5839 9274
rect 5839 9222 5853 9274
rect 5877 9222 5891 9274
rect 5891 9222 5903 9274
rect 5903 9222 5933 9274
rect 5957 9222 5967 9274
rect 5967 9222 6013 9274
rect 5717 9220 5773 9222
rect 5797 9220 5853 9222
rect 5877 9220 5933 9222
rect 5957 9220 6013 9222
rect 5717 8186 5773 8188
rect 5797 8186 5853 8188
rect 5877 8186 5933 8188
rect 5957 8186 6013 8188
rect 5717 8134 5763 8186
rect 5763 8134 5773 8186
rect 5797 8134 5827 8186
rect 5827 8134 5839 8186
rect 5839 8134 5853 8186
rect 5877 8134 5891 8186
rect 5891 8134 5903 8186
rect 5903 8134 5933 8186
rect 5957 8134 5967 8186
rect 5967 8134 6013 8186
rect 5717 8132 5773 8134
rect 5797 8132 5853 8134
rect 5877 8132 5933 8134
rect 5957 8132 6013 8134
rect 5722 7520 5778 7576
rect 5814 7284 5816 7304
rect 5816 7284 5868 7304
rect 5868 7284 5870 7304
rect 5814 7248 5870 7284
rect 5717 7098 5773 7100
rect 5797 7098 5853 7100
rect 5877 7098 5933 7100
rect 5957 7098 6013 7100
rect 5717 7046 5763 7098
rect 5763 7046 5773 7098
rect 5797 7046 5827 7098
rect 5827 7046 5839 7098
rect 5839 7046 5853 7098
rect 5877 7046 5891 7098
rect 5891 7046 5903 7098
rect 5903 7046 5933 7098
rect 5957 7046 5967 7098
rect 5967 7046 6013 7098
rect 5717 7044 5773 7046
rect 5797 7044 5853 7046
rect 5877 7044 5933 7046
rect 5957 7044 6013 7046
rect 4802 3576 4858 3632
rect 5354 5072 5410 5128
rect 5717 6010 5773 6012
rect 5797 6010 5853 6012
rect 5877 6010 5933 6012
rect 5957 6010 6013 6012
rect 5717 5958 5763 6010
rect 5763 5958 5773 6010
rect 5797 5958 5827 6010
rect 5827 5958 5839 6010
rect 5839 5958 5853 6010
rect 5877 5958 5891 6010
rect 5891 5958 5903 6010
rect 5903 5958 5933 6010
rect 5957 5958 5967 6010
rect 5967 5958 6013 6010
rect 5717 5956 5773 5958
rect 5797 5956 5853 5958
rect 5877 5956 5933 5958
rect 5957 5956 6013 5958
rect 5998 5344 6054 5400
rect 6366 9696 6422 9752
rect 7010 12552 7066 12608
rect 7010 11872 7066 11928
rect 6458 8336 6514 8392
rect 6458 6724 6514 6760
rect 6458 6704 6460 6724
rect 6460 6704 6512 6724
rect 6512 6704 6514 6724
rect 5717 4922 5773 4924
rect 5797 4922 5853 4924
rect 5877 4922 5933 4924
rect 5957 4922 6013 4924
rect 5717 4870 5763 4922
rect 5763 4870 5773 4922
rect 5797 4870 5827 4922
rect 5827 4870 5839 4922
rect 5839 4870 5853 4922
rect 5877 4870 5891 4922
rect 5891 4870 5903 4922
rect 5903 4870 5933 4922
rect 5957 4870 5967 4922
rect 5967 4870 6013 4922
rect 5717 4868 5773 4870
rect 5797 4868 5853 4870
rect 5877 4868 5933 4870
rect 5957 4868 6013 4870
rect 6090 4800 6146 4856
rect 5814 4664 5870 4720
rect 5722 3984 5778 4040
rect 5906 4020 5908 4040
rect 5908 4020 5960 4040
rect 5960 4020 5962 4040
rect 5906 3984 5962 4020
rect 5717 3834 5773 3836
rect 5797 3834 5853 3836
rect 5877 3834 5933 3836
rect 5957 3834 6013 3836
rect 5717 3782 5763 3834
rect 5763 3782 5773 3834
rect 5797 3782 5827 3834
rect 5827 3782 5839 3834
rect 5839 3782 5853 3834
rect 5877 3782 5891 3834
rect 5891 3782 5903 3834
rect 5903 3782 5933 3834
rect 5957 3782 5967 3834
rect 5967 3782 6013 3834
rect 5717 3780 5773 3782
rect 5797 3780 5853 3782
rect 5877 3780 5933 3782
rect 5957 3780 6013 3782
rect 4802 2896 4858 2952
rect 5998 3440 6054 3496
rect 5722 3304 5778 3360
rect 5722 3052 5778 3088
rect 5722 3032 5724 3052
rect 5724 3032 5776 3052
rect 5776 3032 5778 3052
rect 5717 2746 5773 2748
rect 5797 2746 5853 2748
rect 5877 2746 5933 2748
rect 5957 2746 6013 2748
rect 5717 2694 5763 2746
rect 5763 2694 5773 2746
rect 5797 2694 5827 2746
rect 5827 2694 5839 2746
rect 5839 2694 5853 2746
rect 5877 2694 5891 2746
rect 5891 2694 5903 2746
rect 5903 2694 5933 2746
rect 5957 2694 5967 2746
rect 5967 2694 6013 2746
rect 5717 2692 5773 2694
rect 5797 2692 5853 2694
rect 5877 2692 5933 2694
rect 5957 2692 6013 2694
rect 6642 4800 6698 4856
rect 7286 12824 7342 12880
rect 7470 13776 7526 13832
rect 8206 17720 8262 17776
rect 8298 15308 8300 15328
rect 8300 15308 8352 15328
rect 8352 15308 8354 15328
rect 7378 12688 7434 12744
rect 7378 12164 7434 12200
rect 7378 12144 7380 12164
rect 7380 12144 7432 12164
rect 7432 12144 7434 12164
rect 7746 12552 7802 12608
rect 7378 10648 7434 10704
rect 7010 8608 7066 8664
rect 7102 8472 7158 8528
rect 8022 13932 8078 13968
rect 8022 13912 8024 13932
rect 8024 13912 8076 13932
rect 8076 13912 8078 13932
rect 8022 12688 8078 12744
rect 8298 15272 8354 15308
rect 8666 16088 8722 16144
rect 8482 15136 8538 15192
rect 8206 13912 8262 13968
rect 8114 11736 8170 11792
rect 8114 11464 8170 11520
rect 6918 6704 6974 6760
rect 7286 6840 7342 6896
rect 7194 6568 7250 6624
rect 6642 2896 6698 2952
rect 6918 2796 6920 2816
rect 6920 2796 6972 2816
rect 6972 2796 6974 2816
rect 6918 2760 6974 2796
rect 7286 3188 7342 3224
rect 7286 3168 7288 3188
rect 7288 3168 7340 3188
rect 7340 3168 7342 3188
rect 7654 8472 7710 8528
rect 7654 7928 7710 7984
rect 7470 4528 7526 4584
rect 8298 11600 8354 11656
rect 8298 11464 8354 11520
rect 8206 10648 8262 10704
rect 8298 9696 8354 9752
rect 8022 7656 8078 7712
rect 8114 7520 8170 7576
rect 8022 6296 8078 6352
rect 7930 3984 7986 4040
rect 7838 3304 7894 3360
rect 8482 11872 8538 11928
rect 8482 11464 8538 11520
rect 9126 15680 9182 15736
rect 8574 4820 8630 4856
rect 8574 4800 8576 4820
rect 8576 4800 8628 4820
rect 8628 4800 8630 4820
rect 9126 9696 9182 9752
rect 8942 7248 8998 7304
rect 10478 26138 10534 26140
rect 10558 26138 10614 26140
rect 10638 26138 10694 26140
rect 10718 26138 10774 26140
rect 10478 26086 10524 26138
rect 10524 26086 10534 26138
rect 10558 26086 10588 26138
rect 10588 26086 10600 26138
rect 10600 26086 10614 26138
rect 10638 26086 10652 26138
rect 10652 26086 10664 26138
rect 10664 26086 10694 26138
rect 10718 26086 10728 26138
rect 10728 26086 10774 26138
rect 10478 26084 10534 26086
rect 10558 26084 10614 26086
rect 10638 26084 10694 26086
rect 10718 26084 10774 26086
rect 10478 25050 10534 25052
rect 10558 25050 10614 25052
rect 10638 25050 10694 25052
rect 10718 25050 10774 25052
rect 10478 24998 10524 25050
rect 10524 24998 10534 25050
rect 10558 24998 10588 25050
rect 10588 24998 10600 25050
rect 10600 24998 10614 25050
rect 10638 24998 10652 25050
rect 10652 24998 10664 25050
rect 10664 24998 10694 25050
rect 10718 24998 10728 25050
rect 10728 24998 10774 25050
rect 10478 24996 10534 24998
rect 10558 24996 10614 24998
rect 10638 24996 10694 24998
rect 10718 24996 10774 24998
rect 10478 23962 10534 23964
rect 10558 23962 10614 23964
rect 10638 23962 10694 23964
rect 10718 23962 10774 23964
rect 10478 23910 10524 23962
rect 10524 23910 10534 23962
rect 10558 23910 10588 23962
rect 10588 23910 10600 23962
rect 10600 23910 10614 23962
rect 10638 23910 10652 23962
rect 10652 23910 10664 23962
rect 10664 23910 10694 23962
rect 10718 23910 10728 23962
rect 10728 23910 10774 23962
rect 10478 23908 10534 23910
rect 10558 23908 10614 23910
rect 10638 23908 10694 23910
rect 10718 23908 10774 23910
rect 10478 22874 10534 22876
rect 10558 22874 10614 22876
rect 10638 22874 10694 22876
rect 10718 22874 10774 22876
rect 10478 22822 10524 22874
rect 10524 22822 10534 22874
rect 10558 22822 10588 22874
rect 10588 22822 10600 22874
rect 10600 22822 10614 22874
rect 10638 22822 10652 22874
rect 10652 22822 10664 22874
rect 10664 22822 10694 22874
rect 10718 22822 10728 22874
rect 10728 22822 10774 22874
rect 10478 22820 10534 22822
rect 10558 22820 10614 22822
rect 10638 22820 10694 22822
rect 10718 22820 10774 22822
rect 10478 21786 10534 21788
rect 10558 21786 10614 21788
rect 10638 21786 10694 21788
rect 10718 21786 10774 21788
rect 10478 21734 10524 21786
rect 10524 21734 10534 21786
rect 10558 21734 10588 21786
rect 10588 21734 10600 21786
rect 10600 21734 10614 21786
rect 10638 21734 10652 21786
rect 10652 21734 10664 21786
rect 10664 21734 10694 21786
rect 10718 21734 10728 21786
rect 10728 21734 10774 21786
rect 10478 21732 10534 21734
rect 10558 21732 10614 21734
rect 10638 21732 10694 21734
rect 10718 21732 10774 21734
rect 9402 12008 9458 12064
rect 9494 11872 9550 11928
rect 10230 19352 10286 19408
rect 9218 6432 9274 6488
rect 9126 5480 9182 5536
rect 10478 20698 10534 20700
rect 10558 20698 10614 20700
rect 10638 20698 10694 20700
rect 10718 20698 10774 20700
rect 10478 20646 10524 20698
rect 10524 20646 10534 20698
rect 10558 20646 10588 20698
rect 10588 20646 10600 20698
rect 10600 20646 10614 20698
rect 10638 20646 10652 20698
rect 10652 20646 10664 20698
rect 10664 20646 10694 20698
rect 10718 20646 10728 20698
rect 10728 20646 10774 20698
rect 10478 20644 10534 20646
rect 10558 20644 10614 20646
rect 10638 20644 10694 20646
rect 10718 20644 10774 20646
rect 10478 19610 10534 19612
rect 10558 19610 10614 19612
rect 10638 19610 10694 19612
rect 10718 19610 10774 19612
rect 10478 19558 10524 19610
rect 10524 19558 10534 19610
rect 10558 19558 10588 19610
rect 10588 19558 10600 19610
rect 10600 19558 10614 19610
rect 10638 19558 10652 19610
rect 10652 19558 10664 19610
rect 10664 19558 10694 19610
rect 10718 19558 10728 19610
rect 10728 19558 10774 19610
rect 10478 19556 10534 19558
rect 10558 19556 10614 19558
rect 10638 19556 10694 19558
rect 10718 19556 10774 19558
rect 10478 18522 10534 18524
rect 10558 18522 10614 18524
rect 10638 18522 10694 18524
rect 10718 18522 10774 18524
rect 10478 18470 10524 18522
rect 10524 18470 10534 18522
rect 10558 18470 10588 18522
rect 10588 18470 10600 18522
rect 10600 18470 10614 18522
rect 10638 18470 10652 18522
rect 10652 18470 10664 18522
rect 10664 18470 10694 18522
rect 10718 18470 10728 18522
rect 10728 18470 10774 18522
rect 10478 18468 10534 18470
rect 10558 18468 10614 18470
rect 10638 18468 10694 18470
rect 10718 18468 10774 18470
rect 10478 17434 10534 17436
rect 10558 17434 10614 17436
rect 10638 17434 10694 17436
rect 10718 17434 10774 17436
rect 10478 17382 10524 17434
rect 10524 17382 10534 17434
rect 10558 17382 10588 17434
rect 10588 17382 10600 17434
rect 10600 17382 10614 17434
rect 10638 17382 10652 17434
rect 10652 17382 10664 17434
rect 10664 17382 10694 17434
rect 10718 17382 10728 17434
rect 10728 17382 10774 17434
rect 10478 17380 10534 17382
rect 10558 17380 10614 17382
rect 10638 17380 10694 17382
rect 10718 17380 10774 17382
rect 10478 16346 10534 16348
rect 10558 16346 10614 16348
rect 10638 16346 10694 16348
rect 10718 16346 10774 16348
rect 10478 16294 10524 16346
rect 10524 16294 10534 16346
rect 10558 16294 10588 16346
rect 10588 16294 10600 16346
rect 10600 16294 10614 16346
rect 10638 16294 10652 16346
rect 10652 16294 10664 16346
rect 10664 16294 10694 16346
rect 10718 16294 10728 16346
rect 10728 16294 10774 16346
rect 10478 16292 10534 16294
rect 10558 16292 10614 16294
rect 10638 16292 10694 16294
rect 10718 16292 10774 16294
rect 10478 15258 10534 15260
rect 10558 15258 10614 15260
rect 10638 15258 10694 15260
rect 10718 15258 10774 15260
rect 10478 15206 10524 15258
rect 10524 15206 10534 15258
rect 10558 15206 10588 15258
rect 10588 15206 10600 15258
rect 10600 15206 10614 15258
rect 10638 15206 10652 15258
rect 10652 15206 10664 15258
rect 10664 15206 10694 15258
rect 10718 15206 10728 15258
rect 10728 15206 10774 15258
rect 10478 15204 10534 15206
rect 10558 15204 10614 15206
rect 10638 15204 10694 15206
rect 10718 15204 10774 15206
rect 10322 14864 10378 14920
rect 11058 19216 11114 19272
rect 11150 16496 11206 16552
rect 11058 15972 11114 16008
rect 11058 15952 11060 15972
rect 11060 15952 11112 15972
rect 11112 15952 11114 15972
rect 11334 15272 11390 15328
rect 10874 14592 10930 14648
rect 10478 14170 10534 14172
rect 10558 14170 10614 14172
rect 10638 14170 10694 14172
rect 10718 14170 10774 14172
rect 10478 14118 10524 14170
rect 10524 14118 10534 14170
rect 10558 14118 10588 14170
rect 10588 14118 10600 14170
rect 10600 14118 10614 14170
rect 10638 14118 10652 14170
rect 10652 14118 10664 14170
rect 10664 14118 10694 14170
rect 10718 14118 10728 14170
rect 10728 14118 10774 14170
rect 10478 14116 10534 14118
rect 10558 14116 10614 14118
rect 10638 14116 10694 14118
rect 10718 14116 10774 14118
rect 9954 12008 10010 12064
rect 9862 11192 9918 11248
rect 9770 10104 9826 10160
rect 9770 9832 9826 9888
rect 9862 9696 9918 9752
rect 9770 9424 9826 9480
rect 9770 8880 9826 8936
rect 9862 7792 9918 7848
rect 9586 6160 9642 6216
rect 9678 5616 9734 5672
rect 9862 6432 9918 6488
rect 7746 1944 7802 2000
rect 10230 12280 10286 12336
rect 10478 13082 10534 13084
rect 10558 13082 10614 13084
rect 10638 13082 10694 13084
rect 10718 13082 10774 13084
rect 10478 13030 10524 13082
rect 10524 13030 10534 13082
rect 10558 13030 10588 13082
rect 10588 13030 10600 13082
rect 10600 13030 10614 13082
rect 10638 13030 10652 13082
rect 10652 13030 10664 13082
rect 10664 13030 10694 13082
rect 10718 13030 10728 13082
rect 10728 13030 10774 13082
rect 10478 13028 10534 13030
rect 10558 13028 10614 13030
rect 10638 13028 10694 13030
rect 10718 13028 10774 13030
rect 10322 12008 10378 12064
rect 10478 11994 10534 11996
rect 10558 11994 10614 11996
rect 10638 11994 10694 11996
rect 10718 11994 10774 11996
rect 10478 11942 10524 11994
rect 10524 11942 10534 11994
rect 10558 11942 10588 11994
rect 10588 11942 10600 11994
rect 10600 11942 10614 11994
rect 10638 11942 10652 11994
rect 10652 11942 10664 11994
rect 10664 11942 10694 11994
rect 10718 11942 10728 11994
rect 10728 11942 10774 11994
rect 10478 11940 10534 11942
rect 10558 11940 10614 11942
rect 10638 11940 10694 11942
rect 10718 11940 10774 11942
rect 10230 11056 10286 11112
rect 10138 8336 10194 8392
rect 10046 6296 10102 6352
rect 10478 10906 10534 10908
rect 10558 10906 10614 10908
rect 10638 10906 10694 10908
rect 10718 10906 10774 10908
rect 10478 10854 10524 10906
rect 10524 10854 10534 10906
rect 10558 10854 10588 10906
rect 10588 10854 10600 10906
rect 10600 10854 10614 10906
rect 10638 10854 10652 10906
rect 10652 10854 10664 10906
rect 10664 10854 10694 10906
rect 10718 10854 10728 10906
rect 10728 10854 10774 10906
rect 10478 10852 10534 10854
rect 10558 10852 10614 10854
rect 10638 10852 10694 10854
rect 10718 10852 10774 10854
rect 10478 9818 10534 9820
rect 10558 9818 10614 9820
rect 10638 9818 10694 9820
rect 10718 9818 10774 9820
rect 10478 9766 10524 9818
rect 10524 9766 10534 9818
rect 10558 9766 10588 9818
rect 10588 9766 10600 9818
rect 10600 9766 10614 9818
rect 10638 9766 10652 9818
rect 10652 9766 10664 9818
rect 10664 9766 10694 9818
rect 10718 9766 10728 9818
rect 10728 9766 10774 9818
rect 10478 9764 10534 9766
rect 10558 9764 10614 9766
rect 10638 9764 10694 9766
rect 10718 9764 10774 9766
rect 10322 9560 10378 9616
rect 10414 9288 10470 9344
rect 10782 9152 10838 9208
rect 10478 8730 10534 8732
rect 10558 8730 10614 8732
rect 10638 8730 10694 8732
rect 10718 8730 10774 8732
rect 10478 8678 10524 8730
rect 10524 8678 10534 8730
rect 10558 8678 10588 8730
rect 10588 8678 10600 8730
rect 10600 8678 10614 8730
rect 10638 8678 10652 8730
rect 10652 8678 10664 8730
rect 10664 8678 10694 8730
rect 10718 8678 10728 8730
rect 10728 8678 10774 8730
rect 10478 8676 10534 8678
rect 10558 8676 10614 8678
rect 10638 8676 10694 8678
rect 10718 8676 10774 8678
rect 10782 8336 10838 8392
rect 10322 7928 10378 7984
rect 10690 7948 10746 7984
rect 10690 7928 10692 7948
rect 10692 7928 10744 7948
rect 10744 7928 10746 7948
rect 10478 7642 10534 7644
rect 10558 7642 10614 7644
rect 10638 7642 10694 7644
rect 10718 7642 10774 7644
rect 10478 7590 10524 7642
rect 10524 7590 10534 7642
rect 10558 7590 10588 7642
rect 10588 7590 10600 7642
rect 10600 7590 10614 7642
rect 10638 7590 10652 7642
rect 10652 7590 10664 7642
rect 10664 7590 10694 7642
rect 10718 7590 10728 7642
rect 10728 7590 10774 7642
rect 10478 7588 10534 7590
rect 10558 7588 10614 7590
rect 10638 7588 10694 7590
rect 10718 7588 10774 7590
rect 10322 7112 10378 7168
rect 11150 11192 11206 11248
rect 11150 10648 11206 10704
rect 11058 9696 11114 9752
rect 11150 8608 11206 8664
rect 10506 7112 10562 7168
rect 10874 6840 10930 6896
rect 10230 5752 10286 5808
rect 10138 4120 10194 4176
rect 10478 6554 10534 6556
rect 10558 6554 10614 6556
rect 10638 6554 10694 6556
rect 10718 6554 10774 6556
rect 10478 6502 10524 6554
rect 10524 6502 10534 6554
rect 10558 6502 10588 6554
rect 10588 6502 10600 6554
rect 10600 6502 10614 6554
rect 10638 6502 10652 6554
rect 10652 6502 10664 6554
rect 10664 6502 10694 6554
rect 10718 6502 10728 6554
rect 10728 6502 10774 6554
rect 10478 6500 10534 6502
rect 10558 6500 10614 6502
rect 10638 6500 10694 6502
rect 10718 6500 10774 6502
rect 10506 6296 10562 6352
rect 11058 6296 11114 6352
rect 10478 5466 10534 5468
rect 10558 5466 10614 5468
rect 10638 5466 10694 5468
rect 10718 5466 10774 5468
rect 10478 5414 10524 5466
rect 10524 5414 10534 5466
rect 10558 5414 10588 5466
rect 10588 5414 10600 5466
rect 10600 5414 10614 5466
rect 10638 5414 10652 5466
rect 10652 5414 10664 5466
rect 10664 5414 10694 5466
rect 10718 5414 10728 5466
rect 10728 5414 10774 5466
rect 10478 5412 10534 5414
rect 10558 5412 10614 5414
rect 10638 5412 10694 5414
rect 10718 5412 10774 5414
rect 10874 4800 10930 4856
rect 12070 15136 12126 15192
rect 11886 15000 11942 15056
rect 12622 20848 12678 20904
rect 12438 15680 12494 15736
rect 11794 14592 11850 14648
rect 12162 15000 12218 15056
rect 11610 13368 11666 13424
rect 11242 8064 11298 8120
rect 11242 7520 11298 7576
rect 11794 11328 11850 11384
rect 12070 12688 12126 12744
rect 11794 10240 11850 10296
rect 11794 9696 11850 9752
rect 11886 9560 11942 9616
rect 12070 10920 12126 10976
rect 12070 9832 12126 9888
rect 11794 9424 11850 9480
rect 11886 9016 11942 9072
rect 11610 8200 11666 8256
rect 11610 5888 11666 5944
rect 10478 4378 10534 4380
rect 10558 4378 10614 4380
rect 10638 4378 10694 4380
rect 10718 4378 10774 4380
rect 10478 4326 10524 4378
rect 10524 4326 10534 4378
rect 10558 4326 10588 4378
rect 10588 4326 10600 4378
rect 10600 4326 10614 4378
rect 10638 4326 10652 4378
rect 10652 4326 10664 4378
rect 10664 4326 10694 4378
rect 10718 4326 10728 4378
rect 10728 4326 10774 4378
rect 10478 4324 10534 4326
rect 10558 4324 10614 4326
rect 10638 4324 10694 4326
rect 10718 4324 10774 4326
rect 10322 4256 10378 4312
rect 10690 4156 10692 4176
rect 10692 4156 10744 4176
rect 10744 4156 10746 4176
rect 10690 4120 10746 4156
rect 10478 3290 10534 3292
rect 10558 3290 10614 3292
rect 10638 3290 10694 3292
rect 10718 3290 10774 3292
rect 10478 3238 10524 3290
rect 10524 3238 10534 3290
rect 10558 3238 10588 3290
rect 10588 3238 10600 3290
rect 10600 3238 10614 3290
rect 10638 3238 10652 3290
rect 10652 3238 10664 3290
rect 10664 3238 10694 3290
rect 10718 3238 10728 3290
rect 10728 3238 10774 3290
rect 10478 3236 10534 3238
rect 10558 3236 10614 3238
rect 10638 3236 10694 3238
rect 10718 3236 10774 3238
rect 11058 3168 11114 3224
rect 11242 3576 11298 3632
rect 12438 14320 12494 14376
rect 12346 14048 12402 14104
rect 15239 26682 15295 26684
rect 15319 26682 15375 26684
rect 15399 26682 15455 26684
rect 15479 26682 15535 26684
rect 15239 26630 15285 26682
rect 15285 26630 15295 26682
rect 15319 26630 15349 26682
rect 15349 26630 15361 26682
rect 15361 26630 15375 26682
rect 15399 26630 15413 26682
rect 15413 26630 15425 26682
rect 15425 26630 15455 26682
rect 15479 26630 15489 26682
rect 15489 26630 15535 26682
rect 15239 26628 15295 26630
rect 15319 26628 15375 26630
rect 15399 26628 15455 26630
rect 15479 26628 15535 26630
rect 13082 24692 13084 24712
rect 13084 24692 13136 24712
rect 13136 24692 13138 24712
rect 13082 24656 13138 24692
rect 12714 15680 12770 15736
rect 12438 12688 12494 12744
rect 12070 7928 12126 7984
rect 12714 12688 12770 12744
rect 12530 9968 12586 10024
rect 13266 15000 13322 15056
rect 13266 14356 13268 14376
rect 13268 14356 13320 14376
rect 13320 14356 13322 14376
rect 13266 14320 13322 14356
rect 13450 19488 13506 19544
rect 13726 20324 13782 20360
rect 13726 20304 13728 20324
rect 13728 20304 13780 20324
rect 13780 20304 13782 20324
rect 13634 19624 13690 19680
rect 13818 16224 13874 16280
rect 13818 15952 13874 16008
rect 13450 14184 13506 14240
rect 13174 13268 13176 13288
rect 13176 13268 13228 13288
rect 13228 13268 13230 13288
rect 13174 13232 13230 13268
rect 13266 12860 13268 12880
rect 13268 12860 13320 12880
rect 13320 12860 13322 12880
rect 13266 12824 13322 12860
rect 13174 12688 13230 12744
rect 13818 14456 13874 14512
rect 14094 19352 14150 19408
rect 13450 12416 13506 12472
rect 13174 11772 13176 11792
rect 13176 11772 13228 11792
rect 13228 11772 13230 11792
rect 13174 11736 13230 11772
rect 12898 10240 12954 10296
rect 12530 9580 12586 9616
rect 12530 9560 12532 9580
rect 12532 9560 12584 9580
rect 12584 9560 12586 9580
rect 12530 9152 12586 9208
rect 12254 7656 12310 7712
rect 12254 4800 12310 4856
rect 12438 6976 12494 7032
rect 12530 6704 12586 6760
rect 12530 6160 12586 6216
rect 12254 3984 12310 4040
rect 9770 2352 9826 2408
rect 10478 2202 10534 2204
rect 10558 2202 10614 2204
rect 10638 2202 10694 2204
rect 10718 2202 10774 2204
rect 10478 2150 10524 2202
rect 10524 2150 10534 2202
rect 10558 2150 10588 2202
rect 10588 2150 10600 2202
rect 10600 2150 10614 2202
rect 10638 2150 10652 2202
rect 10652 2150 10664 2202
rect 10664 2150 10694 2202
rect 10718 2150 10728 2202
rect 10728 2150 10774 2202
rect 10478 2148 10534 2150
rect 10558 2148 10614 2150
rect 10638 2148 10694 2150
rect 10718 2148 10774 2150
rect 13174 9152 13230 9208
rect 13174 8744 13230 8800
rect 13174 6024 13230 6080
rect 13542 11872 13598 11928
rect 14278 19352 14334 19408
rect 14094 13912 14150 13968
rect 15239 25594 15295 25596
rect 15319 25594 15375 25596
rect 15399 25594 15455 25596
rect 15479 25594 15535 25596
rect 15239 25542 15285 25594
rect 15285 25542 15295 25594
rect 15319 25542 15349 25594
rect 15349 25542 15361 25594
rect 15361 25542 15375 25594
rect 15399 25542 15413 25594
rect 15413 25542 15425 25594
rect 15425 25542 15455 25594
rect 15479 25542 15489 25594
rect 15489 25542 15535 25594
rect 15239 25540 15295 25542
rect 15319 25540 15375 25542
rect 15399 25540 15455 25542
rect 15479 25540 15535 25542
rect 15239 24506 15295 24508
rect 15319 24506 15375 24508
rect 15399 24506 15455 24508
rect 15479 24506 15535 24508
rect 15239 24454 15285 24506
rect 15285 24454 15295 24506
rect 15319 24454 15349 24506
rect 15349 24454 15361 24506
rect 15361 24454 15375 24506
rect 15399 24454 15413 24506
rect 15413 24454 15425 24506
rect 15425 24454 15455 24506
rect 15479 24454 15489 24506
rect 15489 24454 15535 24506
rect 15239 24452 15295 24454
rect 15319 24452 15375 24454
rect 15399 24452 15455 24454
rect 15479 24452 15535 24454
rect 14278 15000 14334 15056
rect 14554 15680 14610 15736
rect 13450 10784 13506 10840
rect 13450 9152 13506 9208
rect 13910 9288 13966 9344
rect 13542 6452 13598 6488
rect 13542 6432 13544 6452
rect 13544 6432 13596 6452
rect 13596 6432 13598 6452
rect 13266 5752 13322 5808
rect 13174 4120 13230 4176
rect 13358 4800 13414 4856
rect 13450 3440 13506 3496
rect 13450 3168 13506 3224
rect 14646 13504 14702 13560
rect 14462 12824 14518 12880
rect 14462 12280 14518 12336
rect 14462 10804 14518 10840
rect 14462 10784 14464 10804
rect 14464 10784 14516 10804
rect 14516 10784 14518 10804
rect 14370 9424 14426 9480
rect 15239 23418 15295 23420
rect 15319 23418 15375 23420
rect 15399 23418 15455 23420
rect 15479 23418 15535 23420
rect 15239 23366 15285 23418
rect 15285 23366 15295 23418
rect 15319 23366 15349 23418
rect 15349 23366 15361 23418
rect 15361 23366 15375 23418
rect 15399 23366 15413 23418
rect 15413 23366 15425 23418
rect 15425 23366 15455 23418
rect 15479 23366 15489 23418
rect 15489 23366 15535 23418
rect 15239 23364 15295 23366
rect 15319 23364 15375 23366
rect 15399 23364 15455 23366
rect 15479 23364 15535 23366
rect 15239 22330 15295 22332
rect 15319 22330 15375 22332
rect 15399 22330 15455 22332
rect 15479 22330 15535 22332
rect 15239 22278 15285 22330
rect 15285 22278 15295 22330
rect 15319 22278 15349 22330
rect 15349 22278 15361 22330
rect 15361 22278 15375 22330
rect 15399 22278 15413 22330
rect 15413 22278 15425 22330
rect 15425 22278 15455 22330
rect 15479 22278 15489 22330
rect 15489 22278 15535 22330
rect 15239 22276 15295 22278
rect 15319 22276 15375 22278
rect 15399 22276 15455 22278
rect 15479 22276 15535 22278
rect 15239 21242 15295 21244
rect 15319 21242 15375 21244
rect 15399 21242 15455 21244
rect 15479 21242 15535 21244
rect 15239 21190 15285 21242
rect 15285 21190 15295 21242
rect 15319 21190 15349 21242
rect 15349 21190 15361 21242
rect 15361 21190 15375 21242
rect 15399 21190 15413 21242
rect 15413 21190 15425 21242
rect 15425 21190 15455 21242
rect 15479 21190 15489 21242
rect 15489 21190 15535 21242
rect 15239 21188 15295 21190
rect 15319 21188 15375 21190
rect 15399 21188 15455 21190
rect 15479 21188 15535 21190
rect 15239 20154 15295 20156
rect 15319 20154 15375 20156
rect 15399 20154 15455 20156
rect 15479 20154 15535 20156
rect 15239 20102 15285 20154
rect 15285 20102 15295 20154
rect 15319 20102 15349 20154
rect 15349 20102 15361 20154
rect 15361 20102 15375 20154
rect 15399 20102 15413 20154
rect 15413 20102 15425 20154
rect 15425 20102 15455 20154
rect 15479 20102 15489 20154
rect 15489 20102 15535 20154
rect 15239 20100 15295 20102
rect 15319 20100 15375 20102
rect 15399 20100 15455 20102
rect 15479 20100 15535 20102
rect 15239 19066 15295 19068
rect 15319 19066 15375 19068
rect 15399 19066 15455 19068
rect 15479 19066 15535 19068
rect 15239 19014 15285 19066
rect 15285 19014 15295 19066
rect 15319 19014 15349 19066
rect 15349 19014 15361 19066
rect 15361 19014 15375 19066
rect 15399 19014 15413 19066
rect 15413 19014 15425 19066
rect 15425 19014 15455 19066
rect 15479 19014 15489 19066
rect 15489 19014 15535 19066
rect 15239 19012 15295 19014
rect 15319 19012 15375 19014
rect 15399 19012 15455 19014
rect 15479 19012 15535 19014
rect 15106 18128 15162 18184
rect 15239 17978 15295 17980
rect 15319 17978 15375 17980
rect 15399 17978 15455 17980
rect 15479 17978 15535 17980
rect 15239 17926 15285 17978
rect 15285 17926 15295 17978
rect 15319 17926 15349 17978
rect 15349 17926 15361 17978
rect 15361 17926 15375 17978
rect 15399 17926 15413 17978
rect 15413 17926 15425 17978
rect 15425 17926 15455 17978
rect 15479 17926 15489 17978
rect 15489 17926 15535 17978
rect 15239 17924 15295 17926
rect 15319 17924 15375 17926
rect 15399 17924 15455 17926
rect 15479 17924 15535 17926
rect 15239 16890 15295 16892
rect 15319 16890 15375 16892
rect 15399 16890 15455 16892
rect 15479 16890 15535 16892
rect 15239 16838 15285 16890
rect 15285 16838 15295 16890
rect 15319 16838 15349 16890
rect 15349 16838 15361 16890
rect 15361 16838 15375 16890
rect 15399 16838 15413 16890
rect 15413 16838 15425 16890
rect 15425 16838 15455 16890
rect 15479 16838 15489 16890
rect 15489 16838 15535 16890
rect 15239 16836 15295 16838
rect 15319 16836 15375 16838
rect 15399 16836 15455 16838
rect 15479 16836 15535 16838
rect 15198 15972 15254 16008
rect 15198 15952 15200 15972
rect 15200 15952 15252 15972
rect 15252 15952 15254 15972
rect 15239 15802 15295 15804
rect 15319 15802 15375 15804
rect 15399 15802 15455 15804
rect 15479 15802 15535 15804
rect 15239 15750 15285 15802
rect 15285 15750 15295 15802
rect 15319 15750 15349 15802
rect 15349 15750 15361 15802
rect 15361 15750 15375 15802
rect 15399 15750 15413 15802
rect 15413 15750 15425 15802
rect 15425 15750 15455 15802
rect 15479 15750 15489 15802
rect 15489 15750 15535 15802
rect 15239 15748 15295 15750
rect 15319 15748 15375 15750
rect 15399 15748 15455 15750
rect 15479 15748 15535 15750
rect 16026 19488 16082 19544
rect 15658 18672 15714 18728
rect 15566 15136 15622 15192
rect 15239 14714 15295 14716
rect 15319 14714 15375 14716
rect 15399 14714 15455 14716
rect 15479 14714 15535 14716
rect 15239 14662 15285 14714
rect 15285 14662 15295 14714
rect 15319 14662 15349 14714
rect 15349 14662 15361 14714
rect 15361 14662 15375 14714
rect 15399 14662 15413 14714
rect 15413 14662 15425 14714
rect 15425 14662 15455 14714
rect 15479 14662 15489 14714
rect 15489 14662 15535 14714
rect 15239 14660 15295 14662
rect 15319 14660 15375 14662
rect 15399 14660 15455 14662
rect 15479 14660 15535 14662
rect 15106 14592 15162 14648
rect 15239 13626 15295 13628
rect 15319 13626 15375 13628
rect 15399 13626 15455 13628
rect 15479 13626 15535 13628
rect 15239 13574 15285 13626
rect 15285 13574 15295 13626
rect 15319 13574 15349 13626
rect 15349 13574 15361 13626
rect 15361 13574 15375 13626
rect 15399 13574 15413 13626
rect 15413 13574 15425 13626
rect 15425 13574 15455 13626
rect 15479 13574 15489 13626
rect 15489 13574 15535 13626
rect 15239 13572 15295 13574
rect 15319 13572 15375 13574
rect 15399 13572 15455 13574
rect 15479 13572 15535 13574
rect 15106 12688 15162 12744
rect 15239 12538 15295 12540
rect 15319 12538 15375 12540
rect 15399 12538 15455 12540
rect 15479 12538 15535 12540
rect 15239 12486 15285 12538
rect 15285 12486 15295 12538
rect 15319 12486 15349 12538
rect 15349 12486 15361 12538
rect 15361 12486 15375 12538
rect 15399 12486 15413 12538
rect 15413 12486 15425 12538
rect 15425 12486 15455 12538
rect 15479 12486 15489 12538
rect 15489 12486 15535 12538
rect 15239 12484 15295 12486
rect 15319 12484 15375 12486
rect 15399 12484 15455 12486
rect 15479 12484 15535 12486
rect 15290 12280 15346 12336
rect 16026 14728 16082 14784
rect 16394 19352 16450 19408
rect 17038 25200 17094 25256
rect 16670 14456 16726 14512
rect 16578 13640 16634 13696
rect 16762 13504 16818 13560
rect 16578 13404 16580 13424
rect 16580 13404 16632 13424
rect 16632 13404 16634 13424
rect 16578 13368 16634 13404
rect 15658 11500 15660 11520
rect 15660 11500 15712 11520
rect 15712 11500 15714 11520
rect 15658 11464 15714 11500
rect 15239 11450 15295 11452
rect 15319 11450 15375 11452
rect 15399 11450 15455 11452
rect 15479 11450 15535 11452
rect 15239 11398 15285 11450
rect 15285 11398 15295 11450
rect 15319 11398 15349 11450
rect 15349 11398 15361 11450
rect 15361 11398 15375 11450
rect 15399 11398 15413 11450
rect 15413 11398 15425 11450
rect 15425 11398 15455 11450
rect 15479 11398 15489 11450
rect 15489 11398 15535 11450
rect 15239 11396 15295 11398
rect 15319 11396 15375 11398
rect 15399 11396 15455 11398
rect 15479 11396 15535 11398
rect 15658 11348 15714 11384
rect 15658 11328 15660 11348
rect 15660 11328 15712 11348
rect 15712 11328 15714 11348
rect 15382 11056 15438 11112
rect 15842 12416 15898 12472
rect 16026 12280 16082 12336
rect 15239 10362 15295 10364
rect 15319 10362 15375 10364
rect 15399 10362 15455 10364
rect 15479 10362 15535 10364
rect 15239 10310 15285 10362
rect 15285 10310 15295 10362
rect 15319 10310 15349 10362
rect 15349 10310 15361 10362
rect 15361 10310 15375 10362
rect 15399 10310 15413 10362
rect 15413 10310 15425 10362
rect 15425 10310 15455 10362
rect 15479 10310 15489 10362
rect 15489 10310 15535 10362
rect 15239 10308 15295 10310
rect 15319 10308 15375 10310
rect 15399 10308 15455 10310
rect 15479 10308 15535 10310
rect 15658 10376 15714 10432
rect 15842 10240 15898 10296
rect 15842 9968 15898 10024
rect 14738 9016 14794 9072
rect 14370 8084 14426 8120
rect 14370 8064 14372 8084
rect 14372 8064 14424 8084
rect 14424 8064 14426 8084
rect 14554 6432 14610 6488
rect 15239 9274 15295 9276
rect 15319 9274 15375 9276
rect 15399 9274 15455 9276
rect 15479 9274 15535 9276
rect 15239 9222 15285 9274
rect 15285 9222 15295 9274
rect 15319 9222 15349 9274
rect 15349 9222 15361 9274
rect 15361 9222 15375 9274
rect 15399 9222 15413 9274
rect 15413 9222 15425 9274
rect 15425 9222 15455 9274
rect 15479 9222 15489 9274
rect 15489 9222 15535 9274
rect 15239 9220 15295 9222
rect 15319 9220 15375 9222
rect 15399 9220 15455 9222
rect 15479 9220 15535 9222
rect 15106 9036 15162 9072
rect 15106 9016 15108 9036
rect 15108 9016 15160 9036
rect 15160 9016 15162 9036
rect 15382 9016 15438 9072
rect 16026 10784 16082 10840
rect 16394 12980 16450 13016
rect 16394 12960 16396 12980
rect 16396 12960 16448 12980
rect 16448 12960 16450 12980
rect 16762 13132 16764 13152
rect 16764 13132 16816 13152
rect 16816 13132 16818 13152
rect 16762 13096 16818 13132
rect 16210 10920 16266 10976
rect 16210 10512 16266 10568
rect 16026 9560 16082 9616
rect 16026 9152 16082 9208
rect 15934 8880 15990 8936
rect 15239 8186 15295 8188
rect 15319 8186 15375 8188
rect 15399 8186 15455 8188
rect 15479 8186 15535 8188
rect 15239 8134 15285 8186
rect 15285 8134 15295 8186
rect 15319 8134 15349 8186
rect 15349 8134 15361 8186
rect 15361 8134 15375 8186
rect 15399 8134 15413 8186
rect 15413 8134 15425 8186
rect 15425 8134 15455 8186
rect 15479 8134 15489 8186
rect 15489 8134 15535 8186
rect 15239 8132 15295 8134
rect 15319 8132 15375 8134
rect 15399 8132 15455 8134
rect 15479 8132 15535 8134
rect 15106 8064 15162 8120
rect 14922 7112 14978 7168
rect 15239 7098 15295 7100
rect 15319 7098 15375 7100
rect 15399 7098 15455 7100
rect 15479 7098 15535 7100
rect 15239 7046 15285 7098
rect 15285 7046 15295 7098
rect 15319 7046 15349 7098
rect 15349 7046 15361 7098
rect 15361 7046 15375 7098
rect 15399 7046 15413 7098
rect 15413 7046 15425 7098
rect 15425 7046 15455 7098
rect 15479 7046 15489 7098
rect 15489 7046 15535 7098
rect 15239 7044 15295 7046
rect 15319 7044 15375 7046
rect 15399 7044 15455 7046
rect 15479 7044 15535 7046
rect 15750 7112 15806 7168
rect 15239 6010 15295 6012
rect 15319 6010 15375 6012
rect 15399 6010 15455 6012
rect 15479 6010 15535 6012
rect 15239 5958 15285 6010
rect 15285 5958 15295 6010
rect 15319 5958 15349 6010
rect 15349 5958 15361 6010
rect 15361 5958 15375 6010
rect 15399 5958 15413 6010
rect 15413 5958 15425 6010
rect 15425 5958 15455 6010
rect 15479 5958 15489 6010
rect 15489 5958 15535 6010
rect 15239 5956 15295 5958
rect 15319 5956 15375 5958
rect 15399 5956 15455 5958
rect 15479 5956 15535 5958
rect 14922 5888 14978 5944
rect 14278 5480 14334 5536
rect 13910 3168 13966 3224
rect 14370 4936 14426 4992
rect 14094 3032 14150 3088
rect 14738 5616 14794 5672
rect 15198 5752 15254 5808
rect 14830 5108 14832 5128
rect 14832 5108 14884 5128
rect 14884 5108 14886 5128
rect 14830 5072 14886 5108
rect 15014 5072 15070 5128
rect 15842 6704 15898 6760
rect 15750 6024 15806 6080
rect 15750 5908 15806 5944
rect 15750 5888 15752 5908
rect 15752 5888 15804 5908
rect 15804 5888 15806 5908
rect 15382 5480 15438 5536
rect 15566 5480 15622 5536
rect 15290 5244 15292 5264
rect 15292 5244 15344 5264
rect 15344 5244 15346 5264
rect 15290 5208 15346 5244
rect 15474 5208 15530 5264
rect 15239 4922 15295 4924
rect 15319 4922 15375 4924
rect 15399 4922 15455 4924
rect 15479 4922 15535 4924
rect 15239 4870 15285 4922
rect 15285 4870 15295 4922
rect 15319 4870 15349 4922
rect 15349 4870 15361 4922
rect 15361 4870 15375 4922
rect 15399 4870 15413 4922
rect 15413 4870 15425 4922
rect 15425 4870 15455 4922
rect 15479 4870 15489 4922
rect 15489 4870 15535 4922
rect 15239 4868 15295 4870
rect 15319 4868 15375 4870
rect 15399 4868 15455 4870
rect 15479 4868 15535 4870
rect 14554 4548 14610 4584
rect 14554 4528 14556 4548
rect 14556 4528 14608 4548
rect 14608 4528 14610 4548
rect 15566 4256 15622 4312
rect 15239 3834 15295 3836
rect 15319 3834 15375 3836
rect 15399 3834 15455 3836
rect 15479 3834 15535 3836
rect 15239 3782 15285 3834
rect 15285 3782 15295 3834
rect 15319 3782 15349 3834
rect 15349 3782 15361 3834
rect 15361 3782 15375 3834
rect 15399 3782 15413 3834
rect 15413 3782 15425 3834
rect 15425 3782 15455 3834
rect 15479 3782 15489 3834
rect 15489 3782 15535 3834
rect 15239 3780 15295 3782
rect 15319 3780 15375 3782
rect 15399 3780 15455 3782
rect 15479 3780 15535 3782
rect 13818 2216 13874 2272
rect 13634 2080 13690 2136
rect 13266 1672 13322 1728
rect 15239 2746 15295 2748
rect 15319 2746 15375 2748
rect 15399 2746 15455 2748
rect 15479 2746 15535 2748
rect 15239 2694 15285 2746
rect 15285 2694 15295 2746
rect 15319 2694 15349 2746
rect 15349 2694 15361 2746
rect 15361 2694 15375 2746
rect 15399 2694 15413 2746
rect 15413 2694 15425 2746
rect 15425 2694 15455 2746
rect 15479 2694 15489 2746
rect 15489 2694 15535 2746
rect 15239 2692 15295 2694
rect 15319 2692 15375 2694
rect 15399 2692 15455 2694
rect 15479 2692 15535 2694
rect 20000 26138 20056 26140
rect 20080 26138 20136 26140
rect 20160 26138 20216 26140
rect 20240 26138 20296 26140
rect 20000 26086 20046 26138
rect 20046 26086 20056 26138
rect 20080 26086 20110 26138
rect 20110 26086 20122 26138
rect 20122 26086 20136 26138
rect 20160 26086 20174 26138
rect 20174 26086 20186 26138
rect 20186 26086 20216 26138
rect 20240 26086 20250 26138
rect 20250 26086 20296 26138
rect 20000 26084 20056 26086
rect 20080 26084 20136 26086
rect 20160 26084 20216 26086
rect 20240 26084 20296 26086
rect 17406 18264 17462 18320
rect 17314 15952 17370 16008
rect 17314 15272 17370 15328
rect 16578 11056 16634 11112
rect 16486 9580 16542 9616
rect 16486 9560 16488 9580
rect 16488 9560 16540 9580
rect 16540 9560 16542 9580
rect 16394 6976 16450 7032
rect 17406 15000 17462 15056
rect 17498 14900 17500 14920
rect 17500 14900 17552 14920
rect 17552 14900 17554 14920
rect 17498 14864 17554 14900
rect 17866 18128 17922 18184
rect 17498 12008 17554 12064
rect 17406 11872 17462 11928
rect 17498 11464 17554 11520
rect 16946 11056 17002 11112
rect 16762 7948 16818 7984
rect 16762 7928 16764 7948
rect 16764 7928 16816 7948
rect 16816 7928 16818 7948
rect 17222 9868 17224 9888
rect 17224 9868 17276 9888
rect 17276 9868 17278 9888
rect 17222 9832 17278 9868
rect 17314 8744 17370 8800
rect 17038 8336 17094 8392
rect 16946 7520 17002 7576
rect 17222 8064 17278 8120
rect 17314 7520 17370 7576
rect 16486 6432 16542 6488
rect 16578 6296 16634 6352
rect 16210 5888 16266 5944
rect 16670 5480 16726 5536
rect 16118 5208 16174 5264
rect 16302 4664 16358 4720
rect 16302 4140 16358 4176
rect 16302 4120 16304 4140
rect 16304 4120 16356 4140
rect 16356 4120 16358 4140
rect 15198 2488 15254 2544
rect 17222 7384 17278 7440
rect 17866 14320 17922 14376
rect 17774 12280 17830 12336
rect 17682 11872 17738 11928
rect 17866 12008 17922 12064
rect 17774 11600 17830 11656
rect 17866 11328 17922 11384
rect 17498 8608 17554 8664
rect 17498 7656 17554 7712
rect 17038 3440 17094 3496
rect 17590 6976 17646 7032
rect 17498 6432 17554 6488
rect 17038 2760 17094 2816
rect 17130 2624 17186 2680
rect 17590 6024 17646 6080
rect 17774 9424 17830 9480
rect 17958 6568 18014 6624
rect 17958 3984 18014 4040
rect 18694 20712 18750 20768
rect 20000 25050 20056 25052
rect 20080 25050 20136 25052
rect 20160 25050 20216 25052
rect 20240 25050 20296 25052
rect 20000 24998 20046 25050
rect 20046 24998 20056 25050
rect 20080 24998 20110 25050
rect 20110 24998 20122 25050
rect 20122 24998 20136 25050
rect 20160 24998 20174 25050
rect 20174 24998 20186 25050
rect 20186 24998 20216 25050
rect 20240 24998 20250 25050
rect 20250 24998 20296 25050
rect 20000 24996 20056 24998
rect 20080 24996 20136 24998
rect 20160 24996 20216 24998
rect 20240 24996 20296 24998
rect 19154 20984 19210 21040
rect 20000 23962 20056 23964
rect 20080 23962 20136 23964
rect 20160 23962 20216 23964
rect 20240 23962 20296 23964
rect 20000 23910 20046 23962
rect 20046 23910 20056 23962
rect 20080 23910 20110 23962
rect 20110 23910 20122 23962
rect 20122 23910 20136 23962
rect 20160 23910 20174 23962
rect 20174 23910 20186 23962
rect 20186 23910 20216 23962
rect 20240 23910 20250 23962
rect 20250 23910 20296 23962
rect 20000 23908 20056 23910
rect 20080 23908 20136 23910
rect 20160 23908 20216 23910
rect 20240 23908 20296 23910
rect 20000 22874 20056 22876
rect 20080 22874 20136 22876
rect 20160 22874 20216 22876
rect 20240 22874 20296 22876
rect 20000 22822 20046 22874
rect 20046 22822 20056 22874
rect 20080 22822 20110 22874
rect 20110 22822 20122 22874
rect 20122 22822 20136 22874
rect 20160 22822 20174 22874
rect 20174 22822 20186 22874
rect 20186 22822 20216 22874
rect 20240 22822 20250 22874
rect 20250 22822 20296 22874
rect 20000 22820 20056 22822
rect 20080 22820 20136 22822
rect 20160 22820 20216 22822
rect 20240 22820 20296 22822
rect 19338 19896 19394 19952
rect 18694 16768 18750 16824
rect 18510 14728 18566 14784
rect 18602 14048 18658 14104
rect 18510 12960 18566 13016
rect 18786 13524 18842 13560
rect 18786 13504 18788 13524
rect 18788 13504 18840 13524
rect 18840 13504 18842 13524
rect 18326 4256 18382 4312
rect 18234 3984 18290 4040
rect 18602 10920 18658 10976
rect 19062 12960 19118 13016
rect 18694 9696 18750 9752
rect 19338 19624 19394 19680
rect 19338 17312 19394 17368
rect 19522 16904 19578 16960
rect 19430 14900 19432 14920
rect 19432 14900 19484 14920
rect 19484 14900 19486 14920
rect 19430 14864 19486 14900
rect 20000 21786 20056 21788
rect 20080 21786 20136 21788
rect 20160 21786 20216 21788
rect 20240 21786 20296 21788
rect 20000 21734 20046 21786
rect 20046 21734 20056 21786
rect 20080 21734 20110 21786
rect 20110 21734 20122 21786
rect 20122 21734 20136 21786
rect 20160 21734 20174 21786
rect 20174 21734 20186 21786
rect 20186 21734 20216 21786
rect 20240 21734 20250 21786
rect 20250 21734 20296 21786
rect 20000 21732 20056 21734
rect 20080 21732 20136 21734
rect 20160 21732 20216 21734
rect 20240 21732 20296 21734
rect 20000 20698 20056 20700
rect 20080 20698 20136 20700
rect 20160 20698 20216 20700
rect 20240 20698 20296 20700
rect 20000 20646 20046 20698
rect 20046 20646 20056 20698
rect 20080 20646 20110 20698
rect 20110 20646 20122 20698
rect 20122 20646 20136 20698
rect 20160 20646 20174 20698
rect 20174 20646 20186 20698
rect 20186 20646 20216 20698
rect 20240 20646 20250 20698
rect 20250 20646 20296 20698
rect 20000 20644 20056 20646
rect 20080 20644 20136 20646
rect 20160 20644 20216 20646
rect 20240 20644 20296 20646
rect 19890 19760 19946 19816
rect 20000 19610 20056 19612
rect 20080 19610 20136 19612
rect 20160 19610 20216 19612
rect 20240 19610 20296 19612
rect 20000 19558 20046 19610
rect 20046 19558 20056 19610
rect 20080 19558 20110 19610
rect 20110 19558 20122 19610
rect 20122 19558 20136 19610
rect 20160 19558 20174 19610
rect 20174 19558 20186 19610
rect 20186 19558 20216 19610
rect 20240 19558 20250 19610
rect 20250 19558 20296 19610
rect 20000 19556 20056 19558
rect 20080 19556 20136 19558
rect 20160 19556 20216 19558
rect 20240 19556 20296 19558
rect 19706 15136 19762 15192
rect 20000 18522 20056 18524
rect 20080 18522 20136 18524
rect 20160 18522 20216 18524
rect 20240 18522 20296 18524
rect 20000 18470 20046 18522
rect 20046 18470 20056 18522
rect 20080 18470 20110 18522
rect 20110 18470 20122 18522
rect 20122 18470 20136 18522
rect 20160 18470 20174 18522
rect 20174 18470 20186 18522
rect 20186 18470 20216 18522
rect 20240 18470 20250 18522
rect 20250 18470 20296 18522
rect 20000 18468 20056 18470
rect 20080 18468 20136 18470
rect 20160 18468 20216 18470
rect 20240 18468 20296 18470
rect 20902 23432 20958 23488
rect 21270 20304 21326 20360
rect 20718 19624 20774 19680
rect 20000 17434 20056 17436
rect 20080 17434 20136 17436
rect 20160 17434 20216 17436
rect 20240 17434 20296 17436
rect 20000 17382 20046 17434
rect 20046 17382 20056 17434
rect 20080 17382 20110 17434
rect 20110 17382 20122 17434
rect 20122 17382 20136 17434
rect 20160 17382 20174 17434
rect 20174 17382 20186 17434
rect 20186 17382 20216 17434
rect 20240 17382 20250 17434
rect 20250 17382 20296 17434
rect 20000 17380 20056 17382
rect 20080 17380 20136 17382
rect 20160 17380 20216 17382
rect 20240 17380 20296 17382
rect 20000 16346 20056 16348
rect 20080 16346 20136 16348
rect 20160 16346 20216 16348
rect 20240 16346 20296 16348
rect 20000 16294 20046 16346
rect 20046 16294 20056 16346
rect 20080 16294 20110 16346
rect 20110 16294 20122 16346
rect 20122 16294 20136 16346
rect 20160 16294 20174 16346
rect 20174 16294 20186 16346
rect 20186 16294 20216 16346
rect 20240 16294 20250 16346
rect 20250 16294 20296 16346
rect 20000 16292 20056 16294
rect 20080 16292 20136 16294
rect 20160 16292 20216 16294
rect 20240 16292 20296 16294
rect 20074 16088 20130 16144
rect 20442 16088 20498 16144
rect 20000 15258 20056 15260
rect 20080 15258 20136 15260
rect 20160 15258 20216 15260
rect 20240 15258 20296 15260
rect 20000 15206 20046 15258
rect 20046 15206 20056 15258
rect 20080 15206 20110 15258
rect 20110 15206 20122 15258
rect 20122 15206 20136 15258
rect 20160 15206 20174 15258
rect 20174 15206 20186 15258
rect 20186 15206 20216 15258
rect 20240 15206 20250 15258
rect 20250 15206 20296 15258
rect 20000 15204 20056 15206
rect 20080 15204 20136 15206
rect 20160 15204 20216 15206
rect 20240 15204 20296 15206
rect 19982 15036 19984 15056
rect 19984 15036 20036 15056
rect 20036 15036 20038 15056
rect 19982 15000 20038 15036
rect 20000 14170 20056 14172
rect 20080 14170 20136 14172
rect 20160 14170 20216 14172
rect 20240 14170 20296 14172
rect 20000 14118 20046 14170
rect 20046 14118 20056 14170
rect 20080 14118 20110 14170
rect 20110 14118 20122 14170
rect 20122 14118 20136 14170
rect 20160 14118 20174 14170
rect 20174 14118 20186 14170
rect 20186 14118 20216 14170
rect 20240 14118 20250 14170
rect 20250 14118 20296 14170
rect 20000 14116 20056 14118
rect 20080 14116 20136 14118
rect 20160 14116 20216 14118
rect 20240 14116 20296 14118
rect 19706 13368 19762 13424
rect 19522 9560 19578 9616
rect 19062 9288 19118 9344
rect 18786 7812 18842 7848
rect 18786 7792 18788 7812
rect 18788 7792 18840 7812
rect 18840 7792 18842 7812
rect 19522 9152 19578 9208
rect 19338 8880 19394 8936
rect 19706 8744 19762 8800
rect 20000 13082 20056 13084
rect 20080 13082 20136 13084
rect 20160 13082 20216 13084
rect 20240 13082 20296 13084
rect 20000 13030 20046 13082
rect 20046 13030 20056 13082
rect 20080 13030 20110 13082
rect 20110 13030 20122 13082
rect 20122 13030 20136 13082
rect 20160 13030 20174 13082
rect 20174 13030 20186 13082
rect 20186 13030 20216 13082
rect 20240 13030 20250 13082
rect 20250 13030 20296 13082
rect 20000 13028 20056 13030
rect 20080 13028 20136 13030
rect 20160 13028 20216 13030
rect 20240 13028 20296 13030
rect 20000 11994 20056 11996
rect 20080 11994 20136 11996
rect 20160 11994 20216 11996
rect 20240 11994 20296 11996
rect 20000 11942 20046 11994
rect 20046 11942 20056 11994
rect 20080 11942 20110 11994
rect 20110 11942 20122 11994
rect 20122 11942 20136 11994
rect 20160 11942 20174 11994
rect 20174 11942 20186 11994
rect 20186 11942 20216 11994
rect 20240 11942 20250 11994
rect 20250 11942 20296 11994
rect 20000 11940 20056 11942
rect 20080 11940 20136 11942
rect 20160 11940 20216 11942
rect 20240 11940 20296 11942
rect 20000 10906 20056 10908
rect 20080 10906 20136 10908
rect 20160 10906 20216 10908
rect 20240 10906 20296 10908
rect 20000 10854 20046 10906
rect 20046 10854 20056 10906
rect 20080 10854 20110 10906
rect 20110 10854 20122 10906
rect 20122 10854 20136 10906
rect 20160 10854 20174 10906
rect 20174 10854 20186 10906
rect 20186 10854 20216 10906
rect 20240 10854 20250 10906
rect 20250 10854 20296 10906
rect 20000 10852 20056 10854
rect 20080 10852 20136 10854
rect 20160 10852 20216 10854
rect 20240 10852 20296 10854
rect 20000 9818 20056 9820
rect 20080 9818 20136 9820
rect 20160 9818 20216 9820
rect 20240 9818 20296 9820
rect 20000 9766 20046 9818
rect 20046 9766 20056 9818
rect 20080 9766 20110 9818
rect 20110 9766 20122 9818
rect 20122 9766 20136 9818
rect 20160 9766 20174 9818
rect 20174 9766 20186 9818
rect 20186 9766 20216 9818
rect 20240 9766 20250 9818
rect 20250 9766 20296 9818
rect 20000 9764 20056 9766
rect 20080 9764 20136 9766
rect 20160 9764 20216 9766
rect 20240 9764 20296 9766
rect 19982 9560 20038 9616
rect 20000 8730 20056 8732
rect 20080 8730 20136 8732
rect 20160 8730 20216 8732
rect 20240 8730 20296 8732
rect 20000 8678 20046 8730
rect 20046 8678 20056 8730
rect 20080 8678 20110 8730
rect 20110 8678 20122 8730
rect 20122 8678 20136 8730
rect 20160 8678 20174 8730
rect 20174 8678 20186 8730
rect 20186 8678 20216 8730
rect 20240 8678 20250 8730
rect 20250 8678 20296 8730
rect 20000 8676 20056 8678
rect 20080 8676 20136 8678
rect 20160 8676 20216 8678
rect 20240 8676 20296 8678
rect 20718 10104 20774 10160
rect 19706 7792 19762 7848
rect 19798 6976 19854 7032
rect 20000 7642 20056 7644
rect 20080 7642 20136 7644
rect 20160 7642 20216 7644
rect 20240 7642 20296 7644
rect 20000 7590 20046 7642
rect 20046 7590 20056 7642
rect 20080 7590 20110 7642
rect 20110 7590 20122 7642
rect 20122 7590 20136 7642
rect 20160 7590 20174 7642
rect 20174 7590 20186 7642
rect 20186 7590 20216 7642
rect 20240 7590 20250 7642
rect 20250 7590 20296 7642
rect 20000 7588 20056 7590
rect 20080 7588 20136 7590
rect 20160 7588 20216 7590
rect 20240 7588 20296 7590
rect 20000 6554 20056 6556
rect 20080 6554 20136 6556
rect 20160 6554 20216 6556
rect 20240 6554 20296 6556
rect 20000 6502 20046 6554
rect 20046 6502 20056 6554
rect 20080 6502 20110 6554
rect 20110 6502 20122 6554
rect 20122 6502 20136 6554
rect 20160 6502 20174 6554
rect 20174 6502 20186 6554
rect 20186 6502 20216 6554
rect 20240 6502 20250 6554
rect 20250 6502 20296 6554
rect 20000 6500 20056 6502
rect 20080 6500 20136 6502
rect 20160 6500 20216 6502
rect 20240 6500 20296 6502
rect 19614 5752 19670 5808
rect 19522 4936 19578 4992
rect 18786 4392 18842 4448
rect 19338 4392 19394 4448
rect 19522 4392 19578 4448
rect 19522 4256 19578 4312
rect 20534 7656 20590 7712
rect 20810 6840 20866 6896
rect 20534 6432 20590 6488
rect 20442 6296 20498 6352
rect 20626 6332 20628 6352
rect 20628 6332 20680 6352
rect 20680 6332 20682 6352
rect 20626 6296 20682 6332
rect 20258 5888 20314 5944
rect 20000 5466 20056 5468
rect 20080 5466 20136 5468
rect 20160 5466 20216 5468
rect 20240 5466 20296 5468
rect 20000 5414 20046 5466
rect 20046 5414 20056 5466
rect 20080 5414 20110 5466
rect 20110 5414 20122 5466
rect 20122 5414 20136 5466
rect 20160 5414 20174 5466
rect 20174 5414 20186 5466
rect 20186 5414 20216 5466
rect 20240 5414 20250 5466
rect 20250 5414 20296 5466
rect 20000 5412 20056 5414
rect 20080 5412 20136 5414
rect 20160 5412 20216 5414
rect 20240 5412 20296 5414
rect 20000 4378 20056 4380
rect 20080 4378 20136 4380
rect 20160 4378 20216 4380
rect 20240 4378 20296 4380
rect 20000 4326 20046 4378
rect 20046 4326 20056 4378
rect 20080 4326 20110 4378
rect 20110 4326 20122 4378
rect 20122 4326 20136 4378
rect 20160 4326 20174 4378
rect 20174 4326 20186 4378
rect 20186 4326 20216 4378
rect 20240 4326 20250 4378
rect 20250 4326 20296 4378
rect 20000 4324 20056 4326
rect 20080 4324 20136 4326
rect 20160 4324 20216 4326
rect 20240 4324 20296 4326
rect 20810 6024 20866 6080
rect 20000 3290 20056 3292
rect 20080 3290 20136 3292
rect 20160 3290 20216 3292
rect 20240 3290 20296 3292
rect 20000 3238 20046 3290
rect 20046 3238 20056 3290
rect 20080 3238 20110 3290
rect 20110 3238 20122 3290
rect 20122 3238 20136 3290
rect 20160 3238 20174 3290
rect 20174 3238 20186 3290
rect 20186 3238 20216 3290
rect 20240 3238 20250 3290
rect 20250 3238 20296 3290
rect 20000 3236 20056 3238
rect 20080 3236 20136 3238
rect 20160 3236 20216 3238
rect 20240 3236 20296 3238
rect 18694 2488 18750 2544
rect 19154 2216 19210 2272
rect 19430 2760 19486 2816
rect 21822 20032 21878 20088
rect 21730 19916 21786 19952
rect 21730 19896 21732 19916
rect 21732 19896 21784 19916
rect 21784 19896 21786 19916
rect 21362 15136 21418 15192
rect 21086 9288 21142 9344
rect 20994 9016 21050 9072
rect 20994 8608 21050 8664
rect 20994 8472 21050 8528
rect 22190 19896 22246 19952
rect 22098 19488 22154 19544
rect 22006 12960 22062 13016
rect 22006 12008 22062 12064
rect 21822 11348 21878 11384
rect 21822 11328 21824 11348
rect 21824 11328 21876 11348
rect 21876 11328 21878 11348
rect 21454 8472 21510 8528
rect 21362 8200 21418 8256
rect 21086 5480 21142 5536
rect 20994 5072 21050 5128
rect 20902 2896 20958 2952
rect 21086 3848 21142 3904
rect 20000 2202 20056 2204
rect 20080 2202 20136 2204
rect 20160 2202 20216 2204
rect 20240 2202 20296 2204
rect 20000 2150 20046 2202
rect 20046 2150 20056 2202
rect 20080 2150 20110 2202
rect 20110 2150 20122 2202
rect 20122 2150 20136 2202
rect 20160 2150 20174 2202
rect 20174 2150 20186 2202
rect 20186 2150 20216 2202
rect 20240 2150 20250 2202
rect 20250 2150 20296 2202
rect 20000 2148 20056 2150
rect 20080 2148 20136 2150
rect 20160 2148 20216 2150
rect 20240 2148 20296 2150
rect 21454 7284 21456 7304
rect 21456 7284 21508 7304
rect 21508 7284 21510 7304
rect 21454 7248 21510 7284
rect 21362 4020 21364 4040
rect 21364 4020 21416 4040
rect 21416 4020 21418 4040
rect 21362 3984 21418 4020
rect 21730 9696 21786 9752
rect 22190 11872 22246 11928
rect 21914 8744 21970 8800
rect 22006 6976 22062 7032
rect 21914 5888 21970 5944
rect 21454 3032 21510 3088
rect 22834 19932 22836 19952
rect 22836 19932 22888 19952
rect 22888 19932 22890 19952
rect 22834 19896 22890 19932
rect 22834 19488 22890 19544
rect 22558 15408 22614 15464
rect 23018 13368 23074 13424
rect 22282 9832 22338 9888
rect 22282 9560 22338 9616
rect 22466 11328 22522 11384
rect 22650 10376 22706 10432
rect 22190 8336 22246 8392
rect 22374 8336 22430 8392
rect 22282 7656 22338 7712
rect 22742 9560 22798 9616
rect 22374 6568 22430 6624
rect 22098 5888 22154 5944
rect 22466 6296 22522 6352
rect 22466 6024 22522 6080
rect 22374 5344 22430 5400
rect 22466 5228 22522 5264
rect 22466 5208 22468 5228
rect 22468 5208 22520 5228
rect 22520 5208 22522 5228
rect 22742 6976 22798 7032
rect 23386 18672 23442 18728
rect 23018 11192 23074 11248
rect 22926 11056 22982 11112
rect 23018 5344 23074 5400
rect 21914 2760 21970 2816
rect 23386 15816 23442 15872
rect 23386 15000 23442 15056
rect 24761 26682 24817 26684
rect 24841 26682 24897 26684
rect 24921 26682 24977 26684
rect 25001 26682 25057 26684
rect 24761 26630 24807 26682
rect 24807 26630 24817 26682
rect 24841 26630 24871 26682
rect 24871 26630 24883 26682
rect 24883 26630 24897 26682
rect 24921 26630 24935 26682
rect 24935 26630 24947 26682
rect 24947 26630 24977 26682
rect 25001 26630 25011 26682
rect 25011 26630 25057 26682
rect 24761 26628 24817 26630
rect 24841 26628 24897 26630
rect 24921 26628 24977 26630
rect 25001 26628 25057 26630
rect 24761 25594 24817 25596
rect 24841 25594 24897 25596
rect 24921 25594 24977 25596
rect 25001 25594 25057 25596
rect 24761 25542 24807 25594
rect 24807 25542 24817 25594
rect 24841 25542 24871 25594
rect 24871 25542 24883 25594
rect 24883 25542 24897 25594
rect 24921 25542 24935 25594
rect 24935 25542 24947 25594
rect 24947 25542 24977 25594
rect 25001 25542 25011 25594
rect 25011 25542 25057 25594
rect 24761 25540 24817 25542
rect 24841 25540 24897 25542
rect 24921 25540 24977 25542
rect 25001 25540 25057 25542
rect 24950 24676 25006 24712
rect 24950 24656 24952 24676
rect 24952 24656 25004 24676
rect 25004 24656 25006 24676
rect 24761 24506 24817 24508
rect 24841 24506 24897 24508
rect 24921 24506 24977 24508
rect 25001 24506 25057 24508
rect 24761 24454 24807 24506
rect 24807 24454 24817 24506
rect 24841 24454 24871 24506
rect 24871 24454 24883 24506
rect 24883 24454 24897 24506
rect 24921 24454 24935 24506
rect 24935 24454 24947 24506
rect 24947 24454 24977 24506
rect 25001 24454 25011 24506
rect 25011 24454 25057 24506
rect 24761 24452 24817 24454
rect 24841 24452 24897 24454
rect 24921 24452 24977 24454
rect 25001 24452 25057 24454
rect 23570 20032 23626 20088
rect 23662 17040 23718 17096
rect 24761 23418 24817 23420
rect 24841 23418 24897 23420
rect 24921 23418 24977 23420
rect 25001 23418 25057 23420
rect 24761 23366 24807 23418
rect 24807 23366 24817 23418
rect 24841 23366 24871 23418
rect 24871 23366 24883 23418
rect 24883 23366 24897 23418
rect 24921 23366 24935 23418
rect 24935 23366 24947 23418
rect 24947 23366 24977 23418
rect 25001 23366 25011 23418
rect 25011 23366 25057 23418
rect 24761 23364 24817 23366
rect 24841 23364 24897 23366
rect 24921 23364 24977 23366
rect 25001 23364 25057 23366
rect 24761 22330 24817 22332
rect 24841 22330 24897 22332
rect 24921 22330 24977 22332
rect 25001 22330 25057 22332
rect 24761 22278 24807 22330
rect 24807 22278 24817 22330
rect 24841 22278 24871 22330
rect 24871 22278 24883 22330
rect 24883 22278 24897 22330
rect 24921 22278 24935 22330
rect 24935 22278 24947 22330
rect 24947 22278 24977 22330
rect 25001 22278 25011 22330
rect 25011 22278 25057 22330
rect 24761 22276 24817 22278
rect 24841 22276 24897 22278
rect 24921 22276 24977 22278
rect 25001 22276 25057 22278
rect 24761 21242 24817 21244
rect 24841 21242 24897 21244
rect 24921 21242 24977 21244
rect 25001 21242 25057 21244
rect 24761 21190 24807 21242
rect 24807 21190 24817 21242
rect 24841 21190 24871 21242
rect 24871 21190 24883 21242
rect 24883 21190 24897 21242
rect 24921 21190 24935 21242
rect 24935 21190 24947 21242
rect 24947 21190 24977 21242
rect 25001 21190 25011 21242
rect 25011 21190 25057 21242
rect 24761 21188 24817 21190
rect 24841 21188 24897 21190
rect 24921 21188 24977 21190
rect 25001 21188 25057 21190
rect 24761 20154 24817 20156
rect 24841 20154 24897 20156
rect 24921 20154 24977 20156
rect 25001 20154 25057 20156
rect 24761 20102 24807 20154
rect 24807 20102 24817 20154
rect 24841 20102 24871 20154
rect 24871 20102 24883 20154
rect 24883 20102 24897 20154
rect 24921 20102 24935 20154
rect 24935 20102 24947 20154
rect 24947 20102 24977 20154
rect 25001 20102 25011 20154
rect 25011 20102 25057 20154
rect 24761 20100 24817 20102
rect 24841 20100 24897 20102
rect 24921 20100 24977 20102
rect 25001 20100 25057 20102
rect 24766 19352 24822 19408
rect 24761 19066 24817 19068
rect 24841 19066 24897 19068
rect 24921 19066 24977 19068
rect 25001 19066 25057 19068
rect 24761 19014 24807 19066
rect 24807 19014 24817 19066
rect 24841 19014 24871 19066
rect 24871 19014 24883 19066
rect 24883 19014 24897 19066
rect 24921 19014 24935 19066
rect 24935 19014 24947 19066
rect 24947 19014 24977 19066
rect 25001 19014 25011 19066
rect 25011 19014 25057 19066
rect 24761 19012 24817 19014
rect 24841 19012 24897 19014
rect 24921 19012 24977 19014
rect 25001 19012 25057 19014
rect 24761 17978 24817 17980
rect 24841 17978 24897 17980
rect 24921 17978 24977 17980
rect 25001 17978 25057 17980
rect 24761 17926 24807 17978
rect 24807 17926 24817 17978
rect 24841 17926 24871 17978
rect 24871 17926 24883 17978
rect 24883 17926 24897 17978
rect 24921 17926 24935 17978
rect 24935 17926 24947 17978
rect 24947 17926 24977 17978
rect 25001 17926 25011 17978
rect 25011 17926 25057 17978
rect 24761 17924 24817 17926
rect 24841 17924 24897 17926
rect 24921 17924 24977 17926
rect 25001 17924 25057 17926
rect 24950 17720 25006 17776
rect 24674 17584 24730 17640
rect 23202 11600 23258 11656
rect 23294 8064 23350 8120
rect 24122 14864 24178 14920
rect 23938 12552 23994 12608
rect 23570 11076 23626 11112
rect 23570 11056 23572 11076
rect 23572 11056 23624 11076
rect 23624 11056 23626 11076
rect 23754 7404 23810 7440
rect 23754 7384 23756 7404
rect 23756 7384 23808 7404
rect 23808 7384 23810 7404
rect 23846 7248 23902 7304
rect 23846 4936 23902 4992
rect 24761 16890 24817 16892
rect 24841 16890 24897 16892
rect 24921 16890 24977 16892
rect 25001 16890 25057 16892
rect 24761 16838 24807 16890
rect 24807 16838 24817 16890
rect 24841 16838 24871 16890
rect 24871 16838 24883 16890
rect 24883 16838 24897 16890
rect 24921 16838 24935 16890
rect 24935 16838 24947 16890
rect 24947 16838 24977 16890
rect 25001 16838 25011 16890
rect 25011 16838 25057 16890
rect 24761 16836 24817 16838
rect 24841 16836 24897 16838
rect 24921 16836 24977 16838
rect 25001 16836 25057 16838
rect 26422 22888 26478 22944
rect 25778 20032 25834 20088
rect 25410 18536 25466 18592
rect 25318 17720 25374 17776
rect 24761 15802 24817 15804
rect 24841 15802 24897 15804
rect 24921 15802 24977 15804
rect 25001 15802 25057 15804
rect 24761 15750 24807 15802
rect 24807 15750 24817 15802
rect 24841 15750 24871 15802
rect 24871 15750 24883 15802
rect 24883 15750 24897 15802
rect 24921 15750 24935 15802
rect 24935 15750 24947 15802
rect 24947 15750 24977 15802
rect 25001 15750 25011 15802
rect 25011 15750 25057 15802
rect 24761 15748 24817 15750
rect 24841 15748 24897 15750
rect 24921 15748 24977 15750
rect 25001 15748 25057 15750
rect 24858 15580 24860 15600
rect 24860 15580 24912 15600
rect 24912 15580 24914 15600
rect 24858 15544 24914 15580
rect 25134 14900 25136 14920
rect 25136 14900 25188 14920
rect 25188 14900 25190 14920
rect 25134 14864 25190 14900
rect 24761 14714 24817 14716
rect 24841 14714 24897 14716
rect 24921 14714 24977 14716
rect 25001 14714 25057 14716
rect 24761 14662 24807 14714
rect 24807 14662 24817 14714
rect 24841 14662 24871 14714
rect 24871 14662 24883 14714
rect 24883 14662 24897 14714
rect 24921 14662 24935 14714
rect 24935 14662 24947 14714
rect 24947 14662 24977 14714
rect 25001 14662 25011 14714
rect 25011 14662 25057 14714
rect 24761 14660 24817 14662
rect 24841 14660 24897 14662
rect 24921 14660 24977 14662
rect 25001 14660 25057 14662
rect 24674 14456 24730 14512
rect 24761 13626 24817 13628
rect 24841 13626 24897 13628
rect 24921 13626 24977 13628
rect 25001 13626 25057 13628
rect 24761 13574 24807 13626
rect 24807 13574 24817 13626
rect 24841 13574 24871 13626
rect 24871 13574 24883 13626
rect 24883 13574 24897 13626
rect 24921 13574 24935 13626
rect 24935 13574 24947 13626
rect 24947 13574 24977 13626
rect 25001 13574 25011 13626
rect 25011 13574 25057 13626
rect 24761 13572 24817 13574
rect 24841 13572 24897 13574
rect 24921 13572 24977 13574
rect 25001 13572 25057 13574
rect 24761 12538 24817 12540
rect 24841 12538 24897 12540
rect 24921 12538 24977 12540
rect 25001 12538 25057 12540
rect 24761 12486 24807 12538
rect 24807 12486 24817 12538
rect 24841 12486 24871 12538
rect 24871 12486 24883 12538
rect 24883 12486 24897 12538
rect 24921 12486 24935 12538
rect 24935 12486 24947 12538
rect 24947 12486 24977 12538
rect 25001 12486 25011 12538
rect 25011 12486 25057 12538
rect 24761 12484 24817 12486
rect 24841 12484 24897 12486
rect 24921 12484 24977 12486
rect 25001 12484 25057 12486
rect 24122 6568 24178 6624
rect 23386 3304 23442 3360
rect 24490 9560 24546 9616
rect 24306 6840 24362 6896
rect 24766 11772 24768 11792
rect 24768 11772 24820 11792
rect 24820 11772 24822 11792
rect 24766 11736 24822 11772
rect 24761 11450 24817 11452
rect 24841 11450 24897 11452
rect 24921 11450 24977 11452
rect 25001 11450 25057 11452
rect 24761 11398 24807 11450
rect 24807 11398 24817 11450
rect 24841 11398 24871 11450
rect 24871 11398 24883 11450
rect 24883 11398 24897 11450
rect 24921 11398 24935 11450
rect 24935 11398 24947 11450
rect 24947 11398 24977 11450
rect 25001 11398 25011 11450
rect 25011 11398 25057 11450
rect 24761 11396 24817 11398
rect 24841 11396 24897 11398
rect 24921 11396 24977 11398
rect 25001 11396 25057 11398
rect 24766 10684 24768 10704
rect 24768 10684 24820 10704
rect 24820 10684 24822 10704
rect 24766 10648 24822 10684
rect 24761 10362 24817 10364
rect 24841 10362 24897 10364
rect 24921 10362 24977 10364
rect 25001 10362 25057 10364
rect 24761 10310 24807 10362
rect 24807 10310 24817 10362
rect 24841 10310 24871 10362
rect 24871 10310 24883 10362
rect 24883 10310 24897 10362
rect 24921 10310 24935 10362
rect 24935 10310 24947 10362
rect 24947 10310 24977 10362
rect 25001 10310 25011 10362
rect 25011 10310 25057 10362
rect 24761 10308 24817 10310
rect 24841 10308 24897 10310
rect 24921 10308 24977 10310
rect 25001 10308 25057 10310
rect 25134 10240 25190 10296
rect 25042 9868 25044 9888
rect 25044 9868 25096 9888
rect 25096 9868 25098 9888
rect 25042 9832 25098 9868
rect 25134 9696 25190 9752
rect 24761 9274 24817 9276
rect 24841 9274 24897 9276
rect 24921 9274 24977 9276
rect 25001 9274 25057 9276
rect 24761 9222 24807 9274
rect 24807 9222 24817 9274
rect 24841 9222 24871 9274
rect 24871 9222 24883 9274
rect 24883 9222 24897 9274
rect 24921 9222 24935 9274
rect 24935 9222 24947 9274
rect 24947 9222 24977 9274
rect 25001 9222 25011 9274
rect 25011 9222 25057 9274
rect 24761 9220 24817 9222
rect 24841 9220 24897 9222
rect 24921 9220 24977 9222
rect 25001 9220 25057 9222
rect 24674 8744 24730 8800
rect 24761 8186 24817 8188
rect 24841 8186 24897 8188
rect 24921 8186 24977 8188
rect 25001 8186 25057 8188
rect 24761 8134 24807 8186
rect 24807 8134 24817 8186
rect 24841 8134 24871 8186
rect 24871 8134 24883 8186
rect 24883 8134 24897 8186
rect 24921 8134 24935 8186
rect 24935 8134 24947 8186
rect 24947 8134 24977 8186
rect 25001 8134 25011 8186
rect 25011 8134 25057 8186
rect 24761 8132 24817 8134
rect 24841 8132 24897 8134
rect 24921 8132 24977 8134
rect 25001 8132 25057 8134
rect 24766 7948 24822 7984
rect 24766 7928 24768 7948
rect 24768 7928 24820 7948
rect 24820 7928 24822 7948
rect 25870 19896 25926 19952
rect 26422 19624 26478 19680
rect 26054 18148 26110 18184
rect 26054 18128 26056 18148
rect 26056 18128 26108 18148
rect 26108 18128 26110 18148
rect 25962 17604 26018 17640
rect 25962 17584 25964 17604
rect 25964 17584 26016 17604
rect 26016 17584 26018 17604
rect 27526 24132 27582 24168
rect 27526 24112 27528 24132
rect 27528 24112 27580 24132
rect 27580 24112 27582 24132
rect 27618 21936 27674 21992
rect 26606 17176 26662 17232
rect 26054 17040 26110 17096
rect 26422 16496 26478 16552
rect 25686 15308 25688 15328
rect 25688 15308 25740 15328
rect 25740 15308 25742 15328
rect 25686 15272 25742 15308
rect 25410 11464 25466 11520
rect 25318 11328 25374 11384
rect 25318 11056 25374 11112
rect 25594 12144 25650 12200
rect 25594 11872 25650 11928
rect 25778 11772 25780 11792
rect 25780 11772 25832 11792
rect 25832 11772 25834 11792
rect 25778 11736 25834 11772
rect 25594 11056 25650 11112
rect 25686 10920 25742 10976
rect 25410 10512 25466 10568
rect 25318 10376 25374 10432
rect 25594 10512 25650 10568
rect 25594 10412 25596 10432
rect 25596 10412 25648 10432
rect 25648 10412 25650 10432
rect 25594 10376 25650 10412
rect 25410 9832 25466 9888
rect 26238 11736 26294 11792
rect 26146 11328 26202 11384
rect 25410 9288 25466 9344
rect 25318 9152 25374 9208
rect 25594 8472 25650 8528
rect 25870 10376 25926 10432
rect 25042 7384 25098 7440
rect 25318 7384 25374 7440
rect 25502 7420 25504 7440
rect 25504 7420 25556 7440
rect 25556 7420 25558 7440
rect 25502 7384 25558 7420
rect 24761 7098 24817 7100
rect 24841 7098 24897 7100
rect 24921 7098 24977 7100
rect 25001 7098 25057 7100
rect 24761 7046 24807 7098
rect 24807 7046 24817 7098
rect 24841 7046 24871 7098
rect 24871 7046 24883 7098
rect 24883 7046 24897 7098
rect 24921 7046 24935 7098
rect 24935 7046 24947 7098
rect 24947 7046 24977 7098
rect 25001 7046 25011 7098
rect 25011 7046 25057 7098
rect 24761 7044 24817 7046
rect 24841 7044 24897 7046
rect 24921 7044 24977 7046
rect 25001 7044 25057 7046
rect 25226 7248 25282 7304
rect 25318 7112 25374 7168
rect 25226 6996 25282 7032
rect 25226 6976 25228 6996
rect 25228 6976 25280 6996
rect 25280 6976 25282 6996
rect 25318 6704 25374 6760
rect 24761 6010 24817 6012
rect 24841 6010 24897 6012
rect 24921 6010 24977 6012
rect 25001 6010 25057 6012
rect 24761 5958 24807 6010
rect 24807 5958 24817 6010
rect 24841 5958 24871 6010
rect 24871 5958 24883 6010
rect 24883 5958 24897 6010
rect 24921 5958 24935 6010
rect 24935 5958 24947 6010
rect 24947 5958 24977 6010
rect 25001 5958 25011 6010
rect 25011 5958 25057 6010
rect 24761 5956 24817 5958
rect 24841 5956 24897 5958
rect 24921 5956 24977 5958
rect 25001 5956 25057 5958
rect 24766 5636 24822 5672
rect 24766 5616 24768 5636
rect 24768 5616 24820 5636
rect 24820 5616 24822 5636
rect 25962 9288 26018 9344
rect 25962 9016 26018 9072
rect 29182 26444 29238 26480
rect 29182 26424 29184 26444
rect 29184 26424 29236 26444
rect 29236 26424 29238 26444
rect 26790 13776 26846 13832
rect 26790 12824 26846 12880
rect 26054 7948 26110 7984
rect 26054 7928 26056 7948
rect 26056 7928 26108 7948
rect 26108 7928 26110 7948
rect 25594 5888 25650 5944
rect 26054 7656 26110 7712
rect 27066 17992 27122 18048
rect 27526 17856 27582 17912
rect 29522 26138 29578 26140
rect 29602 26138 29658 26140
rect 29682 26138 29738 26140
rect 29762 26138 29818 26140
rect 29522 26086 29568 26138
rect 29568 26086 29578 26138
rect 29602 26086 29632 26138
rect 29632 26086 29644 26138
rect 29644 26086 29658 26138
rect 29682 26086 29696 26138
rect 29696 26086 29708 26138
rect 29708 26086 29738 26138
rect 29762 26086 29772 26138
rect 29772 26086 29818 26138
rect 29522 26084 29578 26086
rect 29602 26084 29658 26086
rect 29682 26084 29738 26086
rect 29762 26084 29818 26086
rect 28354 19352 28410 19408
rect 27066 16632 27122 16688
rect 26974 12552 27030 12608
rect 26790 10376 26846 10432
rect 25502 5208 25558 5264
rect 25778 4936 25834 4992
rect 24761 4922 24817 4924
rect 24841 4922 24897 4924
rect 24921 4922 24977 4924
rect 25001 4922 25057 4924
rect 24761 4870 24807 4922
rect 24807 4870 24817 4922
rect 24841 4870 24871 4922
rect 24871 4870 24883 4922
rect 24883 4870 24897 4922
rect 24921 4870 24935 4922
rect 24935 4870 24947 4922
rect 24947 4870 24977 4922
rect 25001 4870 25011 4922
rect 25011 4870 25057 4922
rect 24761 4868 24817 4870
rect 24841 4868 24897 4870
rect 24921 4868 24977 4870
rect 25001 4868 25057 4870
rect 25134 3848 25190 3904
rect 24761 3834 24817 3836
rect 24841 3834 24897 3836
rect 24921 3834 24977 3836
rect 25001 3834 25057 3836
rect 24761 3782 24807 3834
rect 24807 3782 24817 3834
rect 24841 3782 24871 3834
rect 24871 3782 24883 3834
rect 24883 3782 24897 3834
rect 24921 3782 24935 3834
rect 24935 3782 24947 3834
rect 24947 3782 24977 3834
rect 25001 3782 25011 3834
rect 25011 3782 25057 3834
rect 24761 3780 24817 3782
rect 24841 3780 24897 3782
rect 24921 3780 24977 3782
rect 25001 3780 25057 3782
rect 26054 3984 26110 4040
rect 26422 7656 26478 7712
rect 26422 5888 26478 5944
rect 26330 4664 26386 4720
rect 26330 4392 26386 4448
rect 25962 3848 26018 3904
rect 26146 3476 26148 3496
rect 26148 3476 26200 3496
rect 26200 3476 26202 3496
rect 26146 3440 26202 3476
rect 24761 2746 24817 2748
rect 24841 2746 24897 2748
rect 24921 2746 24977 2748
rect 25001 2746 25057 2748
rect 24761 2694 24807 2746
rect 24807 2694 24817 2746
rect 24841 2694 24871 2746
rect 24871 2694 24883 2746
rect 24883 2694 24897 2746
rect 24921 2694 24935 2746
rect 24935 2694 24947 2746
rect 24947 2694 24977 2746
rect 25001 2694 25011 2746
rect 25011 2694 25057 2746
rect 24761 2692 24817 2694
rect 24841 2692 24897 2694
rect 24921 2692 24977 2694
rect 25001 2692 25057 2694
rect 25134 2624 25190 2680
rect 25318 2488 25374 2544
rect 26698 6840 26754 6896
rect 27158 9696 27214 9752
rect 27066 7520 27122 7576
rect 26790 5072 26846 5128
rect 26606 3168 26662 3224
rect 27526 11228 27528 11248
rect 27528 11228 27580 11248
rect 27580 11228 27582 11248
rect 27526 11192 27582 11228
rect 27526 10784 27582 10840
rect 27434 10376 27490 10432
rect 27434 10104 27490 10160
rect 27710 9560 27766 9616
rect 27710 7520 27766 7576
rect 28446 17040 28502 17096
rect 29522 25050 29578 25052
rect 29602 25050 29658 25052
rect 29682 25050 29738 25052
rect 29762 25050 29818 25052
rect 29522 24998 29568 25050
rect 29568 24998 29578 25050
rect 29602 24998 29632 25050
rect 29632 24998 29644 25050
rect 29644 24998 29658 25050
rect 29682 24998 29696 25050
rect 29696 24998 29708 25050
rect 29708 24998 29738 25050
rect 29762 24998 29772 25050
rect 29772 24998 29818 25050
rect 29522 24996 29578 24998
rect 29602 24996 29658 24998
rect 29682 24996 29738 24998
rect 29762 24996 29818 24998
rect 29522 23962 29578 23964
rect 29602 23962 29658 23964
rect 29682 23962 29738 23964
rect 29762 23962 29818 23964
rect 29522 23910 29568 23962
rect 29568 23910 29578 23962
rect 29602 23910 29632 23962
rect 29632 23910 29644 23962
rect 29644 23910 29658 23962
rect 29682 23910 29696 23962
rect 29696 23910 29708 23962
rect 29708 23910 29738 23962
rect 29762 23910 29772 23962
rect 29772 23910 29818 23962
rect 29522 23908 29578 23910
rect 29602 23908 29658 23910
rect 29682 23908 29738 23910
rect 29762 23908 29818 23910
rect 29090 18264 29146 18320
rect 28814 16496 28870 16552
rect 28906 15952 28962 16008
rect 27894 13504 27950 13560
rect 27894 11328 27950 11384
rect 27986 11056 28042 11112
rect 27894 9696 27950 9752
rect 27894 9152 27950 9208
rect 28078 8608 28134 8664
rect 27710 6840 27766 6896
rect 27986 8336 28042 8392
rect 28262 9696 28318 9752
rect 28906 15408 28962 15464
rect 29182 15272 29238 15328
rect 28998 13640 29054 13696
rect 29090 13504 29146 13560
rect 29522 22874 29578 22876
rect 29602 22874 29658 22876
rect 29682 22874 29738 22876
rect 29762 22874 29818 22876
rect 29522 22822 29568 22874
rect 29568 22822 29578 22874
rect 29602 22822 29632 22874
rect 29632 22822 29644 22874
rect 29644 22822 29658 22874
rect 29682 22822 29696 22874
rect 29696 22822 29708 22874
rect 29708 22822 29738 22874
rect 29762 22822 29772 22874
rect 29772 22822 29818 22874
rect 29522 22820 29578 22822
rect 29602 22820 29658 22822
rect 29682 22820 29738 22822
rect 29762 22820 29818 22822
rect 29522 21786 29578 21788
rect 29602 21786 29658 21788
rect 29682 21786 29738 21788
rect 29762 21786 29818 21788
rect 29522 21734 29568 21786
rect 29568 21734 29578 21786
rect 29602 21734 29632 21786
rect 29632 21734 29644 21786
rect 29644 21734 29658 21786
rect 29682 21734 29696 21786
rect 29696 21734 29708 21786
rect 29708 21734 29738 21786
rect 29762 21734 29772 21786
rect 29772 21734 29818 21786
rect 29522 21732 29578 21734
rect 29602 21732 29658 21734
rect 29682 21732 29738 21734
rect 29762 21732 29818 21734
rect 29522 20698 29578 20700
rect 29602 20698 29658 20700
rect 29682 20698 29738 20700
rect 29762 20698 29818 20700
rect 29522 20646 29568 20698
rect 29568 20646 29578 20698
rect 29602 20646 29632 20698
rect 29632 20646 29644 20698
rect 29644 20646 29658 20698
rect 29682 20646 29696 20698
rect 29696 20646 29708 20698
rect 29708 20646 29738 20698
rect 29762 20646 29772 20698
rect 29772 20646 29818 20698
rect 29522 20644 29578 20646
rect 29602 20644 29658 20646
rect 29682 20644 29738 20646
rect 29762 20644 29818 20646
rect 29522 19610 29578 19612
rect 29602 19610 29658 19612
rect 29682 19610 29738 19612
rect 29762 19610 29818 19612
rect 29522 19558 29568 19610
rect 29568 19558 29578 19610
rect 29602 19558 29632 19610
rect 29632 19558 29644 19610
rect 29644 19558 29658 19610
rect 29682 19558 29696 19610
rect 29696 19558 29708 19610
rect 29708 19558 29738 19610
rect 29762 19558 29772 19610
rect 29772 19558 29818 19610
rect 29522 19556 29578 19558
rect 29602 19556 29658 19558
rect 29682 19556 29738 19558
rect 29762 19556 29818 19558
rect 29522 18522 29578 18524
rect 29602 18522 29658 18524
rect 29682 18522 29738 18524
rect 29762 18522 29818 18524
rect 29522 18470 29568 18522
rect 29568 18470 29578 18522
rect 29602 18470 29632 18522
rect 29632 18470 29644 18522
rect 29644 18470 29658 18522
rect 29682 18470 29696 18522
rect 29696 18470 29708 18522
rect 29708 18470 29738 18522
rect 29762 18470 29772 18522
rect 29772 18470 29818 18522
rect 29522 18468 29578 18470
rect 29602 18468 29658 18470
rect 29682 18468 29738 18470
rect 29762 18468 29818 18470
rect 29366 17584 29422 17640
rect 29522 17434 29578 17436
rect 29602 17434 29658 17436
rect 29682 17434 29738 17436
rect 29762 17434 29818 17436
rect 29522 17382 29568 17434
rect 29568 17382 29578 17434
rect 29602 17382 29632 17434
rect 29632 17382 29644 17434
rect 29644 17382 29658 17434
rect 29682 17382 29696 17434
rect 29696 17382 29708 17434
rect 29708 17382 29738 17434
rect 29762 17382 29772 17434
rect 29772 17382 29818 17434
rect 29522 17380 29578 17382
rect 29602 17380 29658 17382
rect 29682 17380 29738 17382
rect 29762 17380 29818 17382
rect 29734 17176 29790 17232
rect 30194 20032 30250 20088
rect 29522 16346 29578 16348
rect 29602 16346 29658 16348
rect 29682 16346 29738 16348
rect 29762 16346 29818 16348
rect 29522 16294 29568 16346
rect 29568 16294 29578 16346
rect 29602 16294 29632 16346
rect 29632 16294 29644 16346
rect 29644 16294 29658 16346
rect 29682 16294 29696 16346
rect 29696 16294 29708 16346
rect 29708 16294 29738 16346
rect 29762 16294 29772 16346
rect 29772 16294 29818 16346
rect 29522 16292 29578 16294
rect 29602 16292 29658 16294
rect 29682 16292 29738 16294
rect 29762 16292 29818 16294
rect 30102 17040 30158 17096
rect 29522 15258 29578 15260
rect 29602 15258 29658 15260
rect 29682 15258 29738 15260
rect 29762 15258 29818 15260
rect 29522 15206 29568 15258
rect 29568 15206 29578 15258
rect 29602 15206 29632 15258
rect 29632 15206 29644 15258
rect 29644 15206 29658 15258
rect 29682 15206 29696 15258
rect 29696 15206 29708 15258
rect 29708 15206 29738 15258
rect 29762 15206 29772 15258
rect 29772 15206 29818 15258
rect 29522 15204 29578 15206
rect 29602 15204 29658 15206
rect 29682 15204 29738 15206
rect 29762 15204 29818 15206
rect 29522 14170 29578 14172
rect 29602 14170 29658 14172
rect 29682 14170 29738 14172
rect 29762 14170 29818 14172
rect 29522 14118 29568 14170
rect 29568 14118 29578 14170
rect 29602 14118 29632 14170
rect 29632 14118 29644 14170
rect 29644 14118 29658 14170
rect 29682 14118 29696 14170
rect 29696 14118 29708 14170
rect 29708 14118 29738 14170
rect 29762 14118 29772 14170
rect 29772 14118 29818 14170
rect 29522 14116 29578 14118
rect 29602 14116 29658 14118
rect 29682 14116 29738 14118
rect 29762 14116 29818 14118
rect 29522 13082 29578 13084
rect 29602 13082 29658 13084
rect 29682 13082 29738 13084
rect 29762 13082 29818 13084
rect 29522 13030 29568 13082
rect 29568 13030 29578 13082
rect 29602 13030 29632 13082
rect 29632 13030 29644 13082
rect 29644 13030 29658 13082
rect 29682 13030 29696 13082
rect 29696 13030 29708 13082
rect 29708 13030 29738 13082
rect 29762 13030 29772 13082
rect 29772 13030 29818 13082
rect 29522 13028 29578 13030
rect 29602 13028 29658 13030
rect 29682 13028 29738 13030
rect 29762 13028 29818 13030
rect 29522 11994 29578 11996
rect 29602 11994 29658 11996
rect 29682 11994 29738 11996
rect 29762 11994 29818 11996
rect 29522 11942 29568 11994
rect 29568 11942 29578 11994
rect 29602 11942 29632 11994
rect 29632 11942 29644 11994
rect 29644 11942 29658 11994
rect 29682 11942 29696 11994
rect 29696 11942 29708 11994
rect 29708 11942 29738 11994
rect 29762 11942 29772 11994
rect 29772 11942 29818 11994
rect 29522 11940 29578 11942
rect 29602 11940 29658 11942
rect 29682 11940 29738 11942
rect 29762 11940 29818 11942
rect 28722 11464 28778 11520
rect 29090 10548 29092 10568
rect 29092 10548 29144 10568
rect 29144 10548 29146 10568
rect 29090 10512 29146 10548
rect 29522 10906 29578 10908
rect 29602 10906 29658 10908
rect 29682 10906 29738 10908
rect 29762 10906 29818 10908
rect 29522 10854 29568 10906
rect 29568 10854 29578 10906
rect 29602 10854 29632 10906
rect 29632 10854 29644 10906
rect 29644 10854 29658 10906
rect 29682 10854 29696 10906
rect 29696 10854 29708 10906
rect 29708 10854 29738 10906
rect 29762 10854 29772 10906
rect 29772 10854 29818 10906
rect 29522 10852 29578 10854
rect 29602 10852 29658 10854
rect 29682 10852 29738 10854
rect 29762 10852 29818 10854
rect 29826 10512 29882 10568
rect 29522 9818 29578 9820
rect 29602 9818 29658 9820
rect 29682 9818 29738 9820
rect 29762 9818 29818 9820
rect 29522 9766 29568 9818
rect 29568 9766 29578 9818
rect 29602 9766 29632 9818
rect 29632 9766 29644 9818
rect 29644 9766 29658 9818
rect 29682 9766 29696 9818
rect 29696 9766 29708 9818
rect 29708 9766 29738 9818
rect 29762 9766 29772 9818
rect 29772 9766 29818 9818
rect 29522 9764 29578 9766
rect 29602 9764 29658 9766
rect 29682 9764 29738 9766
rect 29762 9764 29818 9766
rect 28722 9560 28778 9616
rect 28998 9560 29054 9616
rect 28078 7928 28134 7984
rect 27802 5888 27858 5944
rect 27434 5208 27490 5264
rect 27618 5480 27674 5536
rect 27802 5516 27804 5536
rect 27804 5516 27856 5536
rect 27856 5516 27858 5536
rect 27802 5480 27858 5516
rect 27434 3732 27490 3768
rect 27434 3712 27436 3732
rect 27436 3712 27488 3732
rect 27488 3712 27490 3732
rect 27526 3168 27582 3224
rect 27434 2760 27490 2816
rect 28998 9424 29054 9480
rect 28906 8628 28962 8664
rect 28906 8608 28908 8628
rect 28908 8608 28960 8628
rect 28960 8608 28962 8628
rect 28630 8064 28686 8120
rect 28262 5752 28318 5808
rect 28538 5888 28594 5944
rect 28814 8064 28870 8120
rect 29522 8730 29578 8732
rect 29602 8730 29658 8732
rect 29682 8730 29738 8732
rect 29762 8730 29818 8732
rect 29522 8678 29568 8730
rect 29568 8678 29578 8730
rect 29602 8678 29632 8730
rect 29632 8678 29644 8730
rect 29644 8678 29658 8730
rect 29682 8678 29696 8730
rect 29696 8678 29708 8730
rect 29708 8678 29738 8730
rect 29762 8678 29772 8730
rect 29772 8678 29818 8730
rect 29522 8676 29578 8678
rect 29602 8676 29658 8678
rect 29682 8676 29738 8678
rect 29762 8676 29818 8678
rect 29366 8064 29422 8120
rect 29826 8064 29882 8120
rect 28630 5752 28686 5808
rect 28446 5652 28448 5672
rect 28448 5652 28500 5672
rect 28500 5652 28502 5672
rect 28446 5616 28502 5652
rect 28446 5208 28502 5264
rect 28906 7692 28908 7712
rect 28908 7692 28960 7712
rect 28960 7692 28962 7712
rect 28906 7656 28962 7692
rect 29522 7642 29578 7644
rect 29602 7642 29658 7644
rect 29682 7642 29738 7644
rect 29762 7642 29818 7644
rect 29522 7590 29568 7642
rect 29568 7590 29578 7642
rect 29602 7590 29632 7642
rect 29632 7590 29644 7642
rect 29644 7590 29658 7642
rect 29682 7590 29696 7642
rect 29696 7590 29708 7642
rect 29708 7590 29738 7642
rect 29762 7590 29772 7642
rect 29772 7590 29818 7642
rect 29522 7588 29578 7590
rect 29602 7588 29658 7590
rect 29682 7588 29738 7590
rect 29762 7588 29818 7590
rect 29918 7520 29974 7576
rect 29918 7248 29974 7304
rect 30010 6840 30066 6896
rect 29522 6554 29578 6556
rect 29602 6554 29658 6556
rect 29682 6554 29738 6556
rect 29762 6554 29818 6556
rect 29522 6502 29568 6554
rect 29568 6502 29578 6554
rect 29602 6502 29632 6554
rect 29632 6502 29644 6554
rect 29644 6502 29658 6554
rect 29682 6502 29696 6554
rect 29696 6502 29708 6554
rect 29708 6502 29738 6554
rect 29762 6502 29772 6554
rect 29772 6502 29818 6554
rect 29522 6500 29578 6502
rect 29602 6500 29658 6502
rect 29682 6500 29738 6502
rect 29762 6500 29818 6502
rect 31390 22344 31446 22400
rect 30654 19488 30710 19544
rect 30746 19372 30802 19408
rect 30746 19352 30748 19372
rect 30748 19352 30800 19372
rect 30800 19352 30802 19372
rect 30378 16632 30434 16688
rect 30654 18844 30656 18864
rect 30656 18844 30708 18864
rect 30708 18844 30710 18864
rect 30654 18808 30710 18844
rect 30654 18672 30710 18728
rect 30470 15408 30526 15464
rect 30378 11872 30434 11928
rect 30286 10920 30342 10976
rect 30194 9696 30250 9752
rect 30286 9152 30342 9208
rect 30286 8608 30342 8664
rect 30286 7928 30342 7984
rect 30010 6432 30066 6488
rect 28814 4800 28870 4856
rect 29274 5480 29330 5536
rect 29522 5466 29578 5468
rect 29602 5466 29658 5468
rect 29682 5466 29738 5468
rect 29762 5466 29818 5468
rect 29522 5414 29568 5466
rect 29568 5414 29578 5466
rect 29602 5414 29632 5466
rect 29632 5414 29644 5466
rect 29644 5414 29658 5466
rect 29682 5414 29696 5466
rect 29696 5414 29708 5466
rect 29708 5414 29738 5466
rect 29762 5414 29772 5466
rect 29772 5414 29818 5466
rect 29522 5412 29578 5414
rect 29602 5412 29658 5414
rect 29682 5412 29738 5414
rect 29762 5412 29818 5414
rect 29918 5344 29974 5400
rect 29522 4378 29578 4380
rect 29602 4378 29658 4380
rect 29682 4378 29738 4380
rect 29762 4378 29818 4380
rect 29522 4326 29568 4378
rect 29568 4326 29578 4378
rect 29602 4326 29632 4378
rect 29632 4326 29644 4378
rect 29644 4326 29658 4378
rect 29682 4326 29696 4378
rect 29696 4326 29708 4378
rect 29708 4326 29738 4378
rect 29762 4326 29772 4378
rect 29772 4326 29818 4378
rect 29522 4324 29578 4326
rect 29602 4324 29658 4326
rect 29682 4324 29738 4326
rect 29762 4324 29818 4326
rect 30010 3984 30066 4040
rect 29522 3290 29578 3292
rect 29602 3290 29658 3292
rect 29682 3290 29738 3292
rect 29762 3290 29818 3292
rect 29522 3238 29568 3290
rect 29568 3238 29578 3290
rect 29602 3238 29632 3290
rect 29632 3238 29644 3290
rect 29644 3238 29658 3290
rect 29682 3238 29696 3290
rect 29696 3238 29708 3290
rect 29708 3238 29738 3290
rect 29762 3238 29772 3290
rect 29772 3238 29818 3290
rect 29522 3236 29578 3238
rect 29602 3236 29658 3238
rect 29682 3236 29738 3238
rect 29762 3236 29818 3238
rect 32770 22072 32826 22128
rect 32862 21836 32864 21856
rect 32864 21836 32916 21856
rect 32916 21836 32918 21856
rect 32862 21800 32918 21836
rect 32770 20712 32826 20768
rect 31666 17856 31722 17912
rect 32494 17756 32496 17776
rect 32496 17756 32548 17776
rect 32548 17756 32550 17776
rect 32494 17720 32550 17756
rect 31574 17076 31576 17096
rect 31576 17076 31628 17096
rect 31628 17076 31630 17096
rect 31574 17040 31630 17076
rect 31482 16088 31538 16144
rect 31574 15952 31630 16008
rect 30562 8336 30618 8392
rect 30562 7656 30618 7712
rect 30470 6296 30526 6352
rect 30378 5616 30434 5672
rect 30470 5208 30526 5264
rect 29522 2202 29578 2204
rect 29602 2202 29658 2204
rect 29682 2202 29738 2204
rect 29762 2202 29818 2204
rect 29522 2150 29568 2202
rect 29568 2150 29578 2202
rect 29602 2150 29632 2202
rect 29632 2150 29644 2202
rect 29644 2150 29658 2202
rect 29682 2150 29696 2202
rect 29696 2150 29708 2202
rect 29708 2150 29738 2202
rect 29762 2150 29772 2202
rect 29772 2150 29818 2202
rect 29522 2148 29578 2150
rect 29602 2148 29658 2150
rect 29682 2148 29738 2150
rect 29762 2148 29818 2150
rect 30746 10784 30802 10840
rect 30746 10240 30802 10296
rect 30838 9560 30894 9616
rect 31206 11636 31208 11656
rect 31208 11636 31260 11656
rect 31260 11636 31262 11656
rect 31022 9016 31078 9072
rect 31022 8744 31078 8800
rect 30930 7656 30986 7712
rect 31022 6976 31078 7032
rect 30930 6840 30986 6896
rect 30746 4800 30802 4856
rect 31022 5344 31078 5400
rect 31206 11600 31262 11636
rect 31206 11056 31262 11112
rect 31758 12552 31814 12608
rect 31206 8372 31208 8392
rect 31208 8372 31260 8392
rect 31260 8372 31262 8392
rect 31206 8336 31262 8372
rect 31390 9696 31446 9752
rect 32034 12280 32090 12336
rect 31390 9288 31446 9344
rect 31390 9016 31446 9072
rect 31298 8200 31354 8256
rect 31206 6976 31262 7032
rect 31850 9152 31906 9208
rect 31114 5208 31170 5264
rect 31390 3984 31446 4040
rect 31666 4528 31722 4584
rect 31574 3848 31630 3904
rect 32126 8744 32182 8800
rect 33138 17040 33194 17096
rect 32862 13232 32918 13288
rect 32586 10240 32642 10296
rect 33414 17584 33470 17640
rect 33046 13676 33048 13696
rect 33048 13676 33100 13696
rect 33100 13676 33102 13696
rect 33046 13640 33102 13676
rect 33138 12688 33194 12744
rect 33230 12416 33286 12472
rect 32862 9832 32918 9888
rect 32678 7404 32734 7440
rect 32678 7384 32680 7404
rect 32680 7384 32732 7404
rect 32732 7384 32734 7404
rect 33138 11464 33194 11520
rect 33322 11464 33378 11520
rect 33046 8336 33102 8392
rect 32954 8200 33010 8256
rect 32862 6976 32918 7032
rect 32678 6432 32734 6488
rect 32402 4936 32458 4992
rect 31758 2760 31814 2816
rect 32402 3848 32458 3904
rect 32586 6160 32642 6216
rect 33230 10240 33286 10296
rect 33322 9016 33378 9072
rect 33322 5616 33378 5672
rect 32678 3848 32734 3904
rect 34283 26682 34339 26684
rect 34363 26682 34419 26684
rect 34443 26682 34499 26684
rect 34523 26682 34579 26684
rect 34283 26630 34329 26682
rect 34329 26630 34339 26682
rect 34363 26630 34393 26682
rect 34393 26630 34405 26682
rect 34405 26630 34419 26682
rect 34443 26630 34457 26682
rect 34457 26630 34469 26682
rect 34469 26630 34499 26682
rect 34523 26630 34533 26682
rect 34533 26630 34579 26682
rect 34283 26628 34339 26630
rect 34363 26628 34419 26630
rect 34443 26628 34499 26630
rect 34523 26628 34579 26630
rect 34283 25594 34339 25596
rect 34363 25594 34419 25596
rect 34443 25594 34499 25596
rect 34523 25594 34579 25596
rect 34283 25542 34329 25594
rect 34329 25542 34339 25594
rect 34363 25542 34393 25594
rect 34393 25542 34405 25594
rect 34405 25542 34419 25594
rect 34443 25542 34457 25594
rect 34457 25542 34469 25594
rect 34469 25542 34499 25594
rect 34523 25542 34533 25594
rect 34533 25542 34579 25594
rect 34283 25540 34339 25542
rect 34363 25540 34419 25542
rect 34443 25540 34499 25542
rect 34523 25540 34579 25542
rect 34283 24506 34339 24508
rect 34363 24506 34419 24508
rect 34443 24506 34499 24508
rect 34523 24506 34579 24508
rect 34283 24454 34329 24506
rect 34329 24454 34339 24506
rect 34363 24454 34393 24506
rect 34393 24454 34405 24506
rect 34405 24454 34419 24506
rect 34443 24454 34457 24506
rect 34457 24454 34469 24506
rect 34469 24454 34499 24506
rect 34523 24454 34533 24506
rect 34533 24454 34579 24506
rect 34283 24452 34339 24454
rect 34363 24452 34419 24454
rect 34443 24452 34499 24454
rect 34523 24452 34579 24454
rect 34283 23418 34339 23420
rect 34363 23418 34419 23420
rect 34443 23418 34499 23420
rect 34523 23418 34579 23420
rect 34283 23366 34329 23418
rect 34329 23366 34339 23418
rect 34363 23366 34393 23418
rect 34393 23366 34405 23418
rect 34405 23366 34419 23418
rect 34443 23366 34457 23418
rect 34457 23366 34469 23418
rect 34469 23366 34499 23418
rect 34523 23366 34533 23418
rect 34533 23366 34579 23418
rect 34283 23364 34339 23366
rect 34363 23364 34419 23366
rect 34443 23364 34499 23366
rect 34523 23364 34579 23366
rect 33690 19760 33746 19816
rect 33690 15952 33746 16008
rect 34283 22330 34339 22332
rect 34363 22330 34419 22332
rect 34443 22330 34499 22332
rect 34523 22330 34579 22332
rect 34283 22278 34329 22330
rect 34329 22278 34339 22330
rect 34363 22278 34393 22330
rect 34393 22278 34405 22330
rect 34405 22278 34419 22330
rect 34443 22278 34457 22330
rect 34457 22278 34469 22330
rect 34469 22278 34499 22330
rect 34523 22278 34533 22330
rect 34533 22278 34579 22330
rect 34283 22276 34339 22278
rect 34363 22276 34419 22278
rect 34443 22276 34499 22278
rect 34523 22276 34579 22278
rect 34283 21242 34339 21244
rect 34363 21242 34419 21244
rect 34443 21242 34499 21244
rect 34523 21242 34579 21244
rect 34283 21190 34329 21242
rect 34329 21190 34339 21242
rect 34363 21190 34393 21242
rect 34393 21190 34405 21242
rect 34405 21190 34419 21242
rect 34443 21190 34457 21242
rect 34457 21190 34469 21242
rect 34469 21190 34499 21242
rect 34523 21190 34533 21242
rect 34533 21190 34579 21242
rect 34283 21188 34339 21190
rect 34363 21188 34419 21190
rect 34443 21188 34499 21190
rect 34523 21188 34579 21190
rect 34283 20154 34339 20156
rect 34363 20154 34419 20156
rect 34443 20154 34499 20156
rect 34523 20154 34579 20156
rect 34283 20102 34329 20154
rect 34329 20102 34339 20154
rect 34363 20102 34393 20154
rect 34393 20102 34405 20154
rect 34405 20102 34419 20154
rect 34443 20102 34457 20154
rect 34457 20102 34469 20154
rect 34469 20102 34499 20154
rect 34523 20102 34533 20154
rect 34533 20102 34579 20154
rect 34283 20100 34339 20102
rect 34363 20100 34419 20102
rect 34443 20100 34499 20102
rect 34523 20100 34579 20102
rect 34702 19352 34758 19408
rect 34283 19066 34339 19068
rect 34363 19066 34419 19068
rect 34443 19066 34499 19068
rect 34523 19066 34579 19068
rect 34283 19014 34329 19066
rect 34329 19014 34339 19066
rect 34363 19014 34393 19066
rect 34393 19014 34405 19066
rect 34405 19014 34419 19066
rect 34443 19014 34457 19066
rect 34457 19014 34469 19066
rect 34469 19014 34499 19066
rect 34523 19014 34533 19066
rect 34533 19014 34579 19066
rect 34283 19012 34339 19014
rect 34363 19012 34419 19014
rect 34443 19012 34499 19014
rect 34523 19012 34579 19014
rect 33966 13504 34022 13560
rect 34283 17978 34339 17980
rect 34363 17978 34419 17980
rect 34443 17978 34499 17980
rect 34523 17978 34579 17980
rect 34283 17926 34329 17978
rect 34329 17926 34339 17978
rect 34363 17926 34393 17978
rect 34393 17926 34405 17978
rect 34405 17926 34419 17978
rect 34443 17926 34457 17978
rect 34457 17926 34469 17978
rect 34469 17926 34499 17978
rect 34523 17926 34533 17978
rect 34533 17926 34579 17978
rect 34283 17924 34339 17926
rect 34363 17924 34419 17926
rect 34443 17924 34499 17926
rect 34523 17924 34579 17926
rect 34150 17196 34206 17232
rect 34150 17176 34152 17196
rect 34152 17176 34204 17196
rect 34204 17176 34206 17196
rect 34283 16890 34339 16892
rect 34363 16890 34419 16892
rect 34443 16890 34499 16892
rect 34523 16890 34579 16892
rect 34283 16838 34329 16890
rect 34329 16838 34339 16890
rect 34363 16838 34393 16890
rect 34393 16838 34405 16890
rect 34405 16838 34419 16890
rect 34443 16838 34457 16890
rect 34457 16838 34469 16890
rect 34469 16838 34499 16890
rect 34523 16838 34533 16890
rect 34533 16838 34579 16890
rect 34283 16836 34339 16838
rect 34363 16836 34419 16838
rect 34443 16836 34499 16838
rect 34523 16836 34579 16838
rect 34334 15952 34390 16008
rect 34283 15802 34339 15804
rect 34363 15802 34419 15804
rect 34443 15802 34499 15804
rect 34523 15802 34579 15804
rect 34283 15750 34329 15802
rect 34329 15750 34339 15802
rect 34363 15750 34393 15802
rect 34393 15750 34405 15802
rect 34405 15750 34419 15802
rect 34443 15750 34457 15802
rect 34457 15750 34469 15802
rect 34469 15750 34499 15802
rect 34523 15750 34533 15802
rect 34533 15750 34579 15802
rect 34283 15748 34339 15750
rect 34363 15748 34419 15750
rect 34443 15748 34499 15750
rect 34523 15748 34579 15750
rect 34283 14714 34339 14716
rect 34363 14714 34419 14716
rect 34443 14714 34499 14716
rect 34523 14714 34579 14716
rect 34283 14662 34329 14714
rect 34329 14662 34339 14714
rect 34363 14662 34393 14714
rect 34393 14662 34405 14714
rect 34405 14662 34419 14714
rect 34443 14662 34457 14714
rect 34457 14662 34469 14714
rect 34469 14662 34499 14714
rect 34523 14662 34533 14714
rect 34533 14662 34579 14714
rect 34283 14660 34339 14662
rect 34363 14660 34419 14662
rect 34443 14660 34499 14662
rect 34523 14660 34579 14662
rect 34886 16496 34942 16552
rect 34283 13626 34339 13628
rect 34363 13626 34419 13628
rect 34443 13626 34499 13628
rect 34523 13626 34579 13628
rect 34283 13574 34329 13626
rect 34329 13574 34339 13626
rect 34363 13574 34393 13626
rect 34393 13574 34405 13626
rect 34405 13574 34419 13626
rect 34443 13574 34457 13626
rect 34457 13574 34469 13626
rect 34469 13574 34499 13626
rect 34523 13574 34533 13626
rect 34533 13574 34579 13626
rect 34283 13572 34339 13574
rect 34363 13572 34419 13574
rect 34443 13572 34499 13574
rect 34523 13572 34579 13574
rect 33782 12416 33838 12472
rect 33966 11056 34022 11112
rect 34150 12588 34152 12608
rect 34152 12588 34204 12608
rect 34204 12588 34206 12608
rect 34150 12552 34206 12588
rect 34283 12538 34339 12540
rect 34363 12538 34419 12540
rect 34443 12538 34499 12540
rect 34523 12538 34579 12540
rect 34283 12486 34329 12538
rect 34329 12486 34339 12538
rect 34363 12486 34393 12538
rect 34393 12486 34405 12538
rect 34405 12486 34419 12538
rect 34443 12486 34457 12538
rect 34457 12486 34469 12538
rect 34469 12486 34499 12538
rect 34523 12486 34533 12538
rect 34533 12486 34579 12538
rect 34283 12484 34339 12486
rect 34363 12484 34419 12486
rect 34443 12484 34499 12486
rect 34523 12484 34579 12486
rect 37554 26308 37610 26344
rect 37554 26288 37556 26308
rect 37556 26288 37608 26308
rect 37608 26288 37610 26308
rect 35162 15036 35164 15056
rect 35164 15036 35216 15056
rect 35216 15036 35218 15056
rect 35162 15000 35218 15036
rect 34283 11450 34339 11452
rect 34363 11450 34419 11452
rect 34443 11450 34499 11452
rect 34523 11450 34579 11452
rect 34283 11398 34329 11450
rect 34329 11398 34339 11450
rect 34363 11398 34393 11450
rect 34393 11398 34405 11450
rect 34405 11398 34419 11450
rect 34443 11398 34457 11450
rect 34457 11398 34469 11450
rect 34469 11398 34499 11450
rect 34523 11398 34533 11450
rect 34533 11398 34579 11450
rect 34283 11396 34339 11398
rect 34363 11396 34419 11398
rect 34443 11396 34499 11398
rect 34523 11396 34579 11398
rect 33690 9152 33746 9208
rect 33782 8900 33838 8936
rect 33782 8880 33784 8900
rect 33784 8880 33836 8900
rect 33836 8880 33838 8900
rect 33966 10376 34022 10432
rect 34058 10240 34114 10296
rect 33506 8064 33562 8120
rect 33506 6840 33562 6896
rect 33690 8064 33746 8120
rect 33598 5616 33654 5672
rect 33598 5480 33654 5536
rect 33414 3068 33416 3088
rect 33416 3068 33468 3088
rect 33468 3068 33470 3088
rect 33414 3032 33470 3068
rect 33230 2624 33286 2680
rect 34058 9560 34114 9616
rect 34283 10362 34339 10364
rect 34363 10362 34419 10364
rect 34443 10362 34499 10364
rect 34523 10362 34579 10364
rect 34283 10310 34329 10362
rect 34329 10310 34339 10362
rect 34363 10310 34393 10362
rect 34393 10310 34405 10362
rect 34405 10310 34419 10362
rect 34443 10310 34457 10362
rect 34457 10310 34469 10362
rect 34469 10310 34499 10362
rect 34523 10310 34533 10362
rect 34533 10310 34579 10362
rect 34283 10308 34339 10310
rect 34363 10308 34419 10310
rect 34443 10308 34499 10310
rect 34523 10308 34579 10310
rect 34518 9596 34520 9616
rect 34520 9596 34572 9616
rect 34572 9596 34574 9616
rect 34518 9560 34574 9596
rect 34283 9274 34339 9276
rect 34363 9274 34419 9276
rect 34443 9274 34499 9276
rect 34523 9274 34579 9276
rect 34283 9222 34329 9274
rect 34329 9222 34339 9274
rect 34363 9222 34393 9274
rect 34393 9222 34405 9274
rect 34405 9222 34419 9274
rect 34443 9222 34457 9274
rect 34457 9222 34469 9274
rect 34469 9222 34499 9274
rect 34523 9222 34533 9274
rect 34533 9222 34579 9274
rect 34283 9220 34339 9222
rect 34363 9220 34419 9222
rect 34443 9220 34499 9222
rect 34523 9220 34579 9222
rect 34610 8744 34666 8800
rect 34283 8186 34339 8188
rect 34363 8186 34419 8188
rect 34443 8186 34499 8188
rect 34523 8186 34579 8188
rect 34283 8134 34329 8186
rect 34329 8134 34339 8186
rect 34363 8134 34393 8186
rect 34393 8134 34405 8186
rect 34405 8134 34419 8186
rect 34443 8134 34457 8186
rect 34457 8134 34469 8186
rect 34469 8134 34499 8186
rect 34523 8134 34533 8186
rect 34533 8134 34579 8186
rect 34283 8132 34339 8134
rect 34363 8132 34419 8134
rect 34443 8132 34499 8134
rect 34523 8132 34579 8134
rect 34058 6568 34114 6624
rect 33966 5888 34022 5944
rect 33782 4800 33838 4856
rect 34283 7098 34339 7100
rect 34363 7098 34419 7100
rect 34443 7098 34499 7100
rect 34523 7098 34579 7100
rect 34283 7046 34329 7098
rect 34329 7046 34339 7098
rect 34363 7046 34393 7098
rect 34393 7046 34405 7098
rect 34405 7046 34419 7098
rect 34443 7046 34457 7098
rect 34457 7046 34469 7098
rect 34469 7046 34499 7098
rect 34523 7046 34533 7098
rect 34533 7046 34579 7098
rect 34283 7044 34339 7046
rect 34363 7044 34419 7046
rect 34443 7044 34499 7046
rect 34523 7044 34579 7046
rect 34242 6840 34298 6896
rect 34283 6010 34339 6012
rect 34363 6010 34419 6012
rect 34443 6010 34499 6012
rect 34523 6010 34579 6012
rect 34283 5958 34329 6010
rect 34329 5958 34339 6010
rect 34363 5958 34393 6010
rect 34393 5958 34405 6010
rect 34405 5958 34419 6010
rect 34443 5958 34457 6010
rect 34457 5958 34469 6010
rect 34469 5958 34499 6010
rect 34523 5958 34533 6010
rect 34533 5958 34579 6010
rect 34283 5956 34339 5958
rect 34363 5956 34419 5958
rect 34443 5956 34499 5958
rect 34523 5956 34579 5958
rect 34702 8064 34758 8120
rect 34978 11736 35034 11792
rect 34978 8608 35034 8664
rect 35438 15544 35494 15600
rect 35254 9696 35310 9752
rect 35530 10784 35586 10840
rect 35714 9832 35770 9888
rect 35162 7520 35218 7576
rect 34886 6704 34942 6760
rect 34283 4922 34339 4924
rect 34363 4922 34419 4924
rect 34443 4922 34499 4924
rect 34523 4922 34579 4924
rect 34283 4870 34329 4922
rect 34329 4870 34339 4922
rect 34363 4870 34393 4922
rect 34393 4870 34405 4922
rect 34405 4870 34419 4922
rect 34443 4870 34457 4922
rect 34457 4870 34469 4922
rect 34469 4870 34499 4922
rect 34523 4870 34533 4922
rect 34533 4870 34579 4922
rect 34283 4868 34339 4870
rect 34363 4868 34419 4870
rect 34443 4868 34499 4870
rect 34523 4868 34579 4870
rect 34283 3834 34339 3836
rect 34363 3834 34419 3836
rect 34443 3834 34499 3836
rect 34523 3834 34579 3836
rect 34283 3782 34329 3834
rect 34329 3782 34339 3834
rect 34363 3782 34393 3834
rect 34393 3782 34405 3834
rect 34405 3782 34419 3834
rect 34443 3782 34457 3834
rect 34457 3782 34469 3834
rect 34469 3782 34499 3834
rect 34523 3782 34533 3834
rect 34533 3782 34579 3834
rect 34283 3780 34339 3782
rect 34363 3780 34419 3782
rect 34443 3780 34499 3782
rect 34523 3780 34579 3782
rect 35254 6704 35310 6760
rect 35254 6160 35310 6216
rect 35438 4664 35494 4720
rect 34150 2760 34206 2816
rect 34283 2746 34339 2748
rect 34363 2746 34419 2748
rect 34443 2746 34499 2748
rect 34523 2746 34579 2748
rect 34283 2694 34329 2746
rect 34329 2694 34339 2746
rect 34363 2694 34393 2746
rect 34393 2694 34405 2746
rect 34405 2694 34419 2746
rect 34443 2694 34457 2746
rect 34457 2694 34469 2746
rect 34469 2694 34499 2746
rect 34523 2694 34533 2746
rect 34533 2694 34579 2746
rect 34283 2692 34339 2694
rect 34363 2692 34419 2694
rect 34443 2692 34499 2694
rect 34523 2692 34579 2694
rect 34702 1264 34758 1320
rect 36174 9968 36230 10024
rect 36266 7812 36322 7848
rect 36266 7792 36268 7812
rect 36268 7792 36320 7812
rect 36320 7792 36322 7812
rect 36082 7248 36138 7304
rect 35898 6432 35954 6488
rect 36082 6568 36138 6624
rect 36174 6316 36230 6352
rect 36174 6296 36176 6316
rect 36176 6296 36228 6316
rect 36228 6296 36230 6316
rect 36266 4004 36322 4040
rect 36266 3984 36268 4004
rect 36268 3984 36320 4004
rect 36320 3984 36322 4004
rect 37186 19488 37242 19544
rect 36634 14320 36690 14376
rect 36542 9596 36544 9616
rect 36544 9596 36596 9616
rect 36596 9596 36598 9616
rect 36542 9560 36598 9596
rect 37370 14492 37372 14512
rect 37372 14492 37424 14512
rect 37424 14492 37426 14512
rect 37370 14456 37426 14492
rect 37186 12824 37242 12880
rect 37094 11872 37150 11928
rect 36910 8880 36966 8936
rect 36910 6704 36966 6760
rect 36818 5208 36874 5264
rect 36634 3612 36636 3632
rect 36636 3612 36688 3632
rect 36688 3612 36690 3632
rect 36634 3576 36690 3612
rect 36910 5092 36966 5128
rect 36910 5072 36912 5092
rect 36912 5072 36964 5092
rect 36964 5072 36966 5092
rect 37186 7656 37242 7712
rect 39394 27920 39450 27976
rect 39044 26138 39100 26140
rect 39124 26138 39180 26140
rect 39204 26138 39260 26140
rect 39284 26138 39340 26140
rect 39044 26086 39090 26138
rect 39090 26086 39100 26138
rect 39124 26086 39154 26138
rect 39154 26086 39166 26138
rect 39166 26086 39180 26138
rect 39204 26086 39218 26138
rect 39218 26086 39230 26138
rect 39230 26086 39260 26138
rect 39284 26086 39294 26138
rect 39294 26086 39340 26138
rect 39044 26084 39100 26086
rect 39124 26084 39180 26086
rect 39204 26084 39260 26086
rect 39284 26084 39340 26086
rect 39394 25880 39450 25936
rect 39044 25050 39100 25052
rect 39124 25050 39180 25052
rect 39204 25050 39260 25052
rect 39284 25050 39340 25052
rect 39044 24998 39090 25050
rect 39090 24998 39100 25050
rect 39124 24998 39154 25050
rect 39154 24998 39166 25050
rect 39166 24998 39180 25050
rect 39204 24998 39218 25050
rect 39218 24998 39230 25050
rect 39230 24998 39260 25050
rect 39284 24998 39294 25050
rect 39294 24998 39340 25050
rect 39044 24996 39100 24998
rect 39124 24996 39180 24998
rect 39204 24996 39260 24998
rect 39284 24996 39340 24998
rect 39394 24520 39450 24576
rect 39044 23962 39100 23964
rect 39124 23962 39180 23964
rect 39204 23962 39260 23964
rect 39284 23962 39340 23964
rect 39044 23910 39090 23962
rect 39090 23910 39100 23962
rect 39124 23910 39154 23962
rect 39154 23910 39166 23962
rect 39166 23910 39180 23962
rect 39204 23910 39218 23962
rect 39218 23910 39230 23962
rect 39230 23910 39260 23962
rect 39284 23910 39294 23962
rect 39294 23910 39340 23962
rect 39044 23908 39100 23910
rect 39124 23908 39180 23910
rect 39204 23908 39260 23910
rect 39284 23908 39340 23910
rect 39044 22874 39100 22876
rect 39124 22874 39180 22876
rect 39204 22874 39260 22876
rect 39284 22874 39340 22876
rect 39044 22822 39090 22874
rect 39090 22822 39100 22874
rect 39124 22822 39154 22874
rect 39154 22822 39166 22874
rect 39166 22822 39180 22874
rect 39204 22822 39218 22874
rect 39218 22822 39230 22874
rect 39230 22822 39260 22874
rect 39284 22822 39294 22874
rect 39294 22822 39340 22874
rect 39044 22820 39100 22822
rect 39124 22820 39180 22822
rect 39204 22820 39260 22822
rect 39284 22820 39340 22822
rect 39044 21786 39100 21788
rect 39124 21786 39180 21788
rect 39204 21786 39260 21788
rect 39284 21786 39340 21788
rect 39044 21734 39090 21786
rect 39090 21734 39100 21786
rect 39124 21734 39154 21786
rect 39154 21734 39166 21786
rect 39166 21734 39180 21786
rect 39204 21734 39218 21786
rect 39218 21734 39230 21786
rect 39230 21734 39260 21786
rect 39284 21734 39294 21786
rect 39294 21734 39340 21786
rect 39044 21732 39100 21734
rect 39124 21732 39180 21734
rect 39204 21732 39260 21734
rect 39284 21732 39340 21734
rect 39044 20698 39100 20700
rect 39124 20698 39180 20700
rect 39204 20698 39260 20700
rect 39284 20698 39340 20700
rect 39044 20646 39090 20698
rect 39090 20646 39100 20698
rect 39124 20646 39154 20698
rect 39154 20646 39166 20698
rect 39166 20646 39180 20698
rect 39204 20646 39218 20698
rect 39218 20646 39230 20698
rect 39230 20646 39260 20698
rect 39284 20646 39294 20698
rect 39294 20646 39340 20698
rect 39044 20644 39100 20646
rect 39124 20644 39180 20646
rect 39204 20644 39260 20646
rect 39284 20644 39340 20646
rect 39394 20440 39450 20496
rect 38474 19896 38530 19952
rect 39044 19610 39100 19612
rect 39124 19610 39180 19612
rect 39204 19610 39260 19612
rect 39284 19610 39340 19612
rect 39044 19558 39090 19610
rect 39090 19558 39100 19610
rect 39124 19558 39154 19610
rect 39154 19558 39166 19610
rect 39166 19558 39180 19610
rect 39204 19558 39218 19610
rect 39218 19558 39230 19610
rect 39230 19558 39260 19610
rect 39284 19558 39294 19610
rect 39294 19558 39340 19610
rect 39044 19556 39100 19558
rect 39124 19556 39180 19558
rect 39204 19556 39260 19558
rect 39284 19556 39340 19558
rect 39044 18522 39100 18524
rect 39124 18522 39180 18524
rect 39204 18522 39260 18524
rect 39284 18522 39340 18524
rect 39044 18470 39090 18522
rect 39090 18470 39100 18522
rect 39124 18470 39154 18522
rect 39154 18470 39166 18522
rect 39166 18470 39180 18522
rect 39204 18470 39218 18522
rect 39218 18470 39230 18522
rect 39230 18470 39260 18522
rect 39284 18470 39294 18522
rect 39294 18470 39340 18522
rect 39044 18468 39100 18470
rect 39124 18468 39180 18470
rect 39204 18468 39260 18470
rect 39284 18468 39340 18470
rect 39044 17434 39100 17436
rect 39124 17434 39180 17436
rect 39204 17434 39260 17436
rect 39284 17434 39340 17436
rect 39044 17382 39090 17434
rect 39090 17382 39100 17434
rect 39124 17382 39154 17434
rect 39154 17382 39166 17434
rect 39166 17382 39180 17434
rect 39204 17382 39218 17434
rect 39218 17382 39230 17434
rect 39230 17382 39260 17434
rect 39284 17382 39294 17434
rect 39294 17382 39340 17434
rect 39044 17380 39100 17382
rect 39124 17380 39180 17382
rect 39204 17380 39260 17382
rect 39284 17380 39340 17382
rect 37646 10648 37702 10704
rect 37370 8472 37426 8528
rect 36818 2932 36820 2952
rect 36820 2932 36872 2952
rect 36872 2932 36874 2952
rect 36818 2896 36874 2932
rect 35898 1808 35954 1864
rect 37278 1944 37334 2000
rect 37554 8064 37610 8120
rect 38198 10104 38254 10160
rect 37738 8064 37794 8120
rect 37738 7964 37740 7984
rect 37740 7964 37792 7984
rect 37792 7964 37794 7984
rect 37738 7928 37794 7964
rect 38198 8336 38254 8392
rect 37646 4120 37702 4176
rect 38658 17060 38714 17096
rect 38658 17040 38660 17060
rect 38660 17040 38712 17060
rect 38712 17040 38714 17060
rect 39044 16346 39100 16348
rect 39124 16346 39180 16348
rect 39204 16346 39260 16348
rect 39284 16346 39340 16348
rect 39044 16294 39090 16346
rect 39090 16294 39100 16346
rect 39124 16294 39154 16346
rect 39154 16294 39166 16346
rect 39166 16294 39180 16346
rect 39204 16294 39218 16346
rect 39218 16294 39230 16346
rect 39230 16294 39260 16346
rect 39284 16294 39294 16346
rect 39294 16294 39340 16346
rect 39044 16292 39100 16294
rect 39124 16292 39180 16294
rect 39204 16292 39260 16294
rect 39284 16292 39340 16294
rect 39044 15258 39100 15260
rect 39124 15258 39180 15260
rect 39204 15258 39260 15260
rect 39284 15258 39340 15260
rect 39044 15206 39090 15258
rect 39090 15206 39100 15258
rect 39124 15206 39154 15258
rect 39154 15206 39166 15258
rect 39166 15206 39180 15258
rect 39204 15206 39218 15258
rect 39218 15206 39230 15258
rect 39230 15206 39260 15258
rect 39284 15206 39294 15258
rect 39294 15206 39340 15258
rect 39044 15204 39100 15206
rect 39124 15204 39180 15206
rect 39204 15204 39260 15206
rect 39284 15204 39340 15206
rect 38658 15020 38714 15056
rect 38658 15000 38660 15020
rect 38660 15000 38712 15020
rect 38712 15000 38714 15020
rect 39044 14170 39100 14172
rect 39124 14170 39180 14172
rect 39204 14170 39260 14172
rect 39284 14170 39340 14172
rect 39044 14118 39090 14170
rect 39090 14118 39100 14170
rect 39124 14118 39154 14170
rect 39154 14118 39166 14170
rect 39166 14118 39180 14170
rect 39204 14118 39218 14170
rect 39218 14118 39230 14170
rect 39230 14118 39260 14170
rect 39284 14118 39294 14170
rect 39294 14118 39340 14170
rect 39044 14116 39100 14118
rect 39124 14116 39180 14118
rect 39204 14116 39260 14118
rect 39284 14116 39340 14118
rect 39044 13082 39100 13084
rect 39124 13082 39180 13084
rect 39204 13082 39260 13084
rect 39284 13082 39340 13084
rect 39044 13030 39090 13082
rect 39090 13030 39100 13082
rect 39124 13030 39154 13082
rect 39154 13030 39166 13082
rect 39166 13030 39180 13082
rect 39204 13030 39218 13082
rect 39218 13030 39230 13082
rect 39230 13030 39260 13082
rect 39284 13030 39294 13082
rect 39294 13030 39340 13082
rect 39044 13028 39100 13030
rect 39124 13028 39180 13030
rect 39204 13028 39260 13030
rect 39284 13028 39340 13030
rect 39394 12824 39450 12880
rect 39044 11994 39100 11996
rect 39124 11994 39180 11996
rect 39204 11994 39260 11996
rect 39284 11994 39340 11996
rect 39044 11942 39090 11994
rect 39090 11942 39100 11994
rect 39124 11942 39154 11994
rect 39154 11942 39166 11994
rect 39166 11942 39180 11994
rect 39204 11942 39218 11994
rect 39218 11942 39230 11994
rect 39230 11942 39260 11994
rect 39284 11942 39294 11994
rect 39294 11942 39340 11994
rect 39044 11940 39100 11942
rect 39124 11940 39180 11942
rect 39204 11940 39260 11942
rect 39284 11940 39340 11942
rect 39394 11076 39450 11112
rect 39394 11056 39396 11076
rect 39396 11056 39448 11076
rect 39448 11056 39450 11076
rect 39044 10906 39100 10908
rect 39124 10906 39180 10908
rect 39204 10906 39260 10908
rect 39284 10906 39340 10908
rect 39044 10854 39090 10906
rect 39090 10854 39100 10906
rect 39124 10854 39154 10906
rect 39154 10854 39166 10906
rect 39166 10854 39180 10906
rect 39204 10854 39218 10906
rect 39218 10854 39230 10906
rect 39230 10854 39260 10906
rect 39284 10854 39294 10906
rect 39294 10854 39340 10906
rect 39044 10852 39100 10854
rect 39124 10852 39180 10854
rect 39204 10852 39260 10854
rect 39284 10852 39340 10854
rect 39044 9818 39100 9820
rect 39124 9818 39180 9820
rect 39204 9818 39260 9820
rect 39284 9818 39340 9820
rect 39044 9766 39090 9818
rect 39090 9766 39100 9818
rect 39124 9766 39154 9818
rect 39154 9766 39166 9818
rect 39166 9766 39180 9818
rect 39204 9766 39218 9818
rect 39218 9766 39230 9818
rect 39230 9766 39260 9818
rect 39284 9766 39294 9818
rect 39294 9766 39340 9818
rect 39044 9764 39100 9766
rect 39124 9764 39180 9766
rect 39204 9764 39260 9766
rect 39284 9764 39340 9766
rect 39394 9560 39450 9616
rect 39044 8730 39100 8732
rect 39124 8730 39180 8732
rect 39204 8730 39260 8732
rect 39284 8730 39340 8732
rect 39044 8678 39090 8730
rect 39090 8678 39100 8730
rect 39124 8678 39154 8730
rect 39154 8678 39166 8730
rect 39166 8678 39180 8730
rect 39204 8678 39218 8730
rect 39218 8678 39230 8730
rect 39230 8678 39260 8730
rect 39284 8678 39294 8730
rect 39294 8678 39340 8730
rect 39044 8676 39100 8678
rect 39124 8676 39180 8678
rect 39204 8676 39260 8678
rect 39284 8676 39340 8678
rect 39044 7642 39100 7644
rect 39124 7642 39180 7644
rect 39204 7642 39260 7644
rect 39284 7642 39340 7644
rect 39044 7590 39090 7642
rect 39090 7590 39100 7642
rect 39124 7590 39154 7642
rect 39154 7590 39166 7642
rect 39166 7590 39180 7642
rect 39204 7590 39218 7642
rect 39218 7590 39230 7642
rect 39230 7590 39260 7642
rect 39284 7590 39294 7642
rect 39294 7590 39340 7642
rect 39044 7588 39100 7590
rect 39124 7588 39180 7590
rect 39204 7588 39260 7590
rect 39284 7588 39340 7590
rect 38658 7384 38714 7440
rect 38474 2372 38530 2408
rect 38474 2352 38476 2372
rect 38476 2352 38528 2372
rect 38528 2352 38530 2372
rect 38198 1672 38254 1728
rect 39044 6554 39100 6556
rect 39124 6554 39180 6556
rect 39204 6554 39260 6556
rect 39284 6554 39340 6556
rect 39044 6502 39090 6554
rect 39090 6502 39100 6554
rect 39124 6502 39154 6554
rect 39154 6502 39166 6554
rect 39166 6502 39180 6554
rect 39204 6502 39218 6554
rect 39218 6502 39230 6554
rect 39230 6502 39260 6554
rect 39284 6502 39294 6554
rect 39294 6502 39340 6554
rect 39044 6500 39100 6502
rect 39124 6500 39180 6502
rect 39204 6500 39260 6502
rect 39284 6500 39340 6502
rect 39044 5466 39100 5468
rect 39124 5466 39180 5468
rect 39204 5466 39260 5468
rect 39284 5466 39340 5468
rect 39044 5414 39090 5466
rect 39090 5414 39100 5466
rect 39124 5414 39154 5466
rect 39154 5414 39166 5466
rect 39166 5414 39180 5466
rect 39204 5414 39218 5466
rect 39218 5414 39230 5466
rect 39230 5414 39260 5466
rect 39284 5414 39294 5466
rect 39294 5414 39340 5466
rect 39044 5412 39100 5414
rect 39124 5412 39180 5414
rect 39204 5412 39260 5414
rect 39284 5412 39340 5414
rect 39044 4378 39100 4380
rect 39124 4378 39180 4380
rect 39204 4378 39260 4380
rect 39284 4378 39340 4380
rect 39044 4326 39090 4378
rect 39090 4326 39100 4378
rect 39124 4326 39154 4378
rect 39154 4326 39166 4378
rect 39166 4326 39180 4378
rect 39204 4326 39218 4378
rect 39218 4326 39230 4378
rect 39230 4326 39260 4378
rect 39284 4326 39294 4378
rect 39294 4326 39340 4378
rect 39044 4324 39100 4326
rect 39124 4324 39180 4326
rect 39204 4324 39260 4326
rect 39284 4324 39340 4326
rect 38658 3460 38714 3496
rect 38658 3440 38660 3460
rect 38660 3440 38712 3460
rect 38712 3440 38714 3460
rect 39044 3290 39100 3292
rect 39124 3290 39180 3292
rect 39204 3290 39260 3292
rect 39284 3290 39340 3292
rect 39044 3238 39090 3290
rect 39090 3238 39100 3290
rect 39124 3238 39154 3290
rect 39154 3238 39166 3290
rect 39166 3238 39180 3290
rect 39204 3238 39218 3290
rect 39218 3238 39230 3290
rect 39230 3238 39260 3290
rect 39284 3238 39294 3290
rect 39294 3238 39340 3290
rect 39044 3236 39100 3238
rect 39124 3236 39180 3238
rect 39204 3236 39260 3238
rect 39284 3236 39340 3238
rect 39044 2202 39100 2204
rect 39124 2202 39180 2204
rect 39204 2202 39260 2204
rect 39284 2202 39340 2204
rect 39044 2150 39090 2202
rect 39090 2150 39100 2202
rect 39124 2150 39154 2202
rect 39154 2150 39166 2202
rect 39166 2150 39180 2202
rect 39204 2150 39218 2202
rect 39218 2150 39230 2202
rect 39230 2150 39260 2202
rect 39284 2150 39294 2202
rect 39294 2150 39340 2202
rect 39044 2148 39100 2150
rect 39124 2148 39180 2150
rect 39204 2148 39260 2150
rect 39284 2148 39340 2150
rect 38658 1944 38714 2000
rect 39394 40 39450 96
<< metal3 >>
rect 0 27978 800 28008
rect 1025 27978 1091 27981
rect 0 27976 1091 27978
rect 0 27920 1030 27976
rect 1086 27920 1091 27976
rect 0 27918 1091 27920
rect 0 27888 800 27918
rect 1025 27915 1091 27918
rect 39389 27978 39455 27981
rect 39566 27978 40366 28008
rect 39389 27976 40366 27978
rect 39389 27920 39394 27976
rect 39450 27920 40366 27976
rect 39389 27918 40366 27920
rect 39389 27915 39455 27918
rect 39566 27888 40366 27918
rect 5707 26688 6023 26689
rect 5707 26624 5713 26688
rect 5777 26624 5793 26688
rect 5857 26624 5873 26688
rect 5937 26624 5953 26688
rect 6017 26624 6023 26688
rect 5707 26623 6023 26624
rect 15229 26688 15545 26689
rect 15229 26624 15235 26688
rect 15299 26624 15315 26688
rect 15379 26624 15395 26688
rect 15459 26624 15475 26688
rect 15539 26624 15545 26688
rect 15229 26623 15545 26624
rect 24751 26688 25067 26689
rect 24751 26624 24757 26688
rect 24821 26624 24837 26688
rect 24901 26624 24917 26688
rect 24981 26624 24997 26688
rect 25061 26624 25067 26688
rect 24751 26623 25067 26624
rect 34273 26688 34589 26689
rect 34273 26624 34279 26688
rect 34343 26624 34359 26688
rect 34423 26624 34439 26688
rect 34503 26624 34519 26688
rect 34583 26624 34589 26688
rect 34273 26623 34589 26624
rect 12014 26420 12020 26484
rect 12084 26482 12090 26484
rect 29177 26482 29243 26485
rect 12084 26480 29243 26482
rect 12084 26424 29182 26480
rect 29238 26424 29243 26480
rect 12084 26422 29243 26424
rect 12084 26420 12090 26422
rect 29177 26419 29243 26422
rect 3049 26346 3115 26349
rect 6310 26346 6316 26348
rect 3049 26344 6316 26346
rect 3049 26288 3054 26344
rect 3110 26288 6316 26344
rect 3049 26286 6316 26288
rect 3049 26283 3115 26286
rect 6310 26284 6316 26286
rect 6380 26284 6386 26348
rect 7925 26346 7991 26349
rect 14774 26346 14780 26348
rect 7925 26344 14780 26346
rect 7925 26288 7930 26344
rect 7986 26288 14780 26344
rect 7925 26286 14780 26288
rect 7925 26283 7991 26286
rect 14774 26284 14780 26286
rect 14844 26284 14850 26348
rect 18638 26284 18644 26348
rect 18708 26346 18714 26348
rect 37549 26346 37615 26349
rect 18708 26344 37615 26346
rect 18708 26288 37554 26344
rect 37610 26288 37615 26344
rect 18708 26286 37615 26288
rect 18708 26284 18714 26286
rect 37549 26283 37615 26286
rect 10468 26144 10784 26145
rect 10468 26080 10474 26144
rect 10538 26080 10554 26144
rect 10618 26080 10634 26144
rect 10698 26080 10714 26144
rect 10778 26080 10784 26144
rect 10468 26079 10784 26080
rect 19990 26144 20306 26145
rect 19990 26080 19996 26144
rect 20060 26080 20076 26144
rect 20140 26080 20156 26144
rect 20220 26080 20236 26144
rect 20300 26080 20306 26144
rect 19990 26079 20306 26080
rect 29512 26144 29828 26145
rect 29512 26080 29518 26144
rect 29582 26080 29598 26144
rect 29662 26080 29678 26144
rect 29742 26080 29758 26144
rect 29822 26080 29828 26144
rect 29512 26079 29828 26080
rect 39034 26144 39350 26145
rect 39034 26080 39040 26144
rect 39104 26080 39120 26144
rect 39184 26080 39200 26144
rect 39264 26080 39280 26144
rect 39344 26080 39350 26144
rect 39034 26079 39350 26080
rect 0 25938 800 25968
rect 933 25938 999 25941
rect 0 25936 999 25938
rect 0 25880 938 25936
rect 994 25880 999 25936
rect 0 25878 999 25880
rect 0 25848 800 25878
rect 933 25875 999 25878
rect 39389 25938 39455 25941
rect 39566 25938 40366 25968
rect 39389 25936 40366 25938
rect 39389 25880 39394 25936
rect 39450 25880 40366 25936
rect 39389 25878 40366 25880
rect 39389 25875 39455 25878
rect 39566 25848 40366 25878
rect 5707 25600 6023 25601
rect 5707 25536 5713 25600
rect 5777 25536 5793 25600
rect 5857 25536 5873 25600
rect 5937 25536 5953 25600
rect 6017 25536 6023 25600
rect 5707 25535 6023 25536
rect 15229 25600 15545 25601
rect 15229 25536 15235 25600
rect 15299 25536 15315 25600
rect 15379 25536 15395 25600
rect 15459 25536 15475 25600
rect 15539 25536 15545 25600
rect 15229 25535 15545 25536
rect 24751 25600 25067 25601
rect 24751 25536 24757 25600
rect 24821 25536 24837 25600
rect 24901 25536 24917 25600
rect 24981 25536 24997 25600
rect 25061 25536 25067 25600
rect 24751 25535 25067 25536
rect 34273 25600 34589 25601
rect 34273 25536 34279 25600
rect 34343 25536 34359 25600
rect 34423 25536 34439 25600
rect 34503 25536 34519 25600
rect 34583 25536 34589 25600
rect 34273 25535 34589 25536
rect 17033 25258 17099 25261
rect 23974 25258 23980 25260
rect 17033 25256 23980 25258
rect 17033 25200 17038 25256
rect 17094 25200 23980 25256
rect 17033 25198 23980 25200
rect 17033 25195 17099 25198
rect 23974 25196 23980 25198
rect 24044 25196 24050 25260
rect 10468 25056 10784 25057
rect 10468 24992 10474 25056
rect 10538 24992 10554 25056
rect 10618 24992 10634 25056
rect 10698 24992 10714 25056
rect 10778 24992 10784 25056
rect 10468 24991 10784 24992
rect 19990 25056 20306 25057
rect 19990 24992 19996 25056
rect 20060 24992 20076 25056
rect 20140 24992 20156 25056
rect 20220 24992 20236 25056
rect 20300 24992 20306 25056
rect 19990 24991 20306 24992
rect 29512 25056 29828 25057
rect 29512 24992 29518 25056
rect 29582 24992 29598 25056
rect 29662 24992 29678 25056
rect 29742 24992 29758 25056
rect 29822 24992 29828 25056
rect 29512 24991 29828 24992
rect 39034 25056 39350 25057
rect 39034 24992 39040 25056
rect 39104 24992 39120 25056
rect 39184 24992 39200 25056
rect 39264 24992 39280 25056
rect 39344 24992 39350 25056
rect 39034 24991 39350 24992
rect 13077 24716 13143 24717
rect 13077 24714 13124 24716
rect 13032 24712 13124 24714
rect 13032 24656 13082 24712
rect 13032 24654 13124 24656
rect 13077 24652 13124 24654
rect 13188 24652 13194 24716
rect 16614 24652 16620 24716
rect 16684 24714 16690 24716
rect 24945 24714 25011 24717
rect 16684 24712 25011 24714
rect 16684 24656 24950 24712
rect 25006 24656 25011 24712
rect 16684 24654 25011 24656
rect 16684 24652 16690 24654
rect 13077 24651 13143 24652
rect 24945 24651 25011 24654
rect 39389 24578 39455 24581
rect 39566 24578 40366 24608
rect 39389 24576 40366 24578
rect 39389 24520 39394 24576
rect 39450 24520 40366 24576
rect 39389 24518 40366 24520
rect 39389 24515 39455 24518
rect 5707 24512 6023 24513
rect 5707 24448 5713 24512
rect 5777 24448 5793 24512
rect 5857 24448 5873 24512
rect 5937 24448 5953 24512
rect 6017 24448 6023 24512
rect 5707 24447 6023 24448
rect 15229 24512 15545 24513
rect 15229 24448 15235 24512
rect 15299 24448 15315 24512
rect 15379 24448 15395 24512
rect 15459 24448 15475 24512
rect 15539 24448 15545 24512
rect 15229 24447 15545 24448
rect 24751 24512 25067 24513
rect 24751 24448 24757 24512
rect 24821 24448 24837 24512
rect 24901 24448 24917 24512
rect 24981 24448 24997 24512
rect 25061 24448 25067 24512
rect 24751 24447 25067 24448
rect 34273 24512 34589 24513
rect 34273 24448 34279 24512
rect 34343 24448 34359 24512
rect 34423 24448 34439 24512
rect 34503 24448 34519 24512
rect 34583 24448 34589 24512
rect 39566 24488 40366 24518
rect 34273 24447 34589 24448
rect 17166 24108 17172 24172
rect 17236 24170 17242 24172
rect 27521 24170 27587 24173
rect 17236 24168 27587 24170
rect 17236 24112 27526 24168
rect 27582 24112 27587 24168
rect 17236 24110 27587 24112
rect 17236 24108 17242 24110
rect 27521 24107 27587 24110
rect 10468 23968 10784 23969
rect 0 23898 800 23928
rect 10468 23904 10474 23968
rect 10538 23904 10554 23968
rect 10618 23904 10634 23968
rect 10698 23904 10714 23968
rect 10778 23904 10784 23968
rect 10468 23903 10784 23904
rect 19990 23968 20306 23969
rect 19990 23904 19996 23968
rect 20060 23904 20076 23968
rect 20140 23904 20156 23968
rect 20220 23904 20236 23968
rect 20300 23904 20306 23968
rect 19990 23903 20306 23904
rect 29512 23968 29828 23969
rect 29512 23904 29518 23968
rect 29582 23904 29598 23968
rect 29662 23904 29678 23968
rect 29742 23904 29758 23968
rect 29822 23904 29828 23968
rect 29512 23903 29828 23904
rect 39034 23968 39350 23969
rect 39034 23904 39040 23968
rect 39104 23904 39120 23968
rect 39184 23904 39200 23968
rect 39264 23904 39280 23968
rect 39344 23904 39350 23968
rect 39034 23903 39350 23904
rect 933 23898 999 23901
rect 0 23896 999 23898
rect 0 23840 938 23896
rect 994 23840 999 23896
rect 0 23838 999 23840
rect 0 23808 800 23838
rect 933 23835 999 23838
rect 18822 23428 18828 23492
rect 18892 23490 18898 23492
rect 20897 23490 20963 23493
rect 18892 23488 20963 23490
rect 18892 23432 20902 23488
rect 20958 23432 20963 23488
rect 18892 23430 20963 23432
rect 18892 23428 18898 23430
rect 20897 23427 20963 23430
rect 5707 23424 6023 23425
rect 5707 23360 5713 23424
rect 5777 23360 5793 23424
rect 5857 23360 5873 23424
rect 5937 23360 5953 23424
rect 6017 23360 6023 23424
rect 5707 23359 6023 23360
rect 15229 23424 15545 23425
rect 15229 23360 15235 23424
rect 15299 23360 15315 23424
rect 15379 23360 15395 23424
rect 15459 23360 15475 23424
rect 15539 23360 15545 23424
rect 15229 23359 15545 23360
rect 24751 23424 25067 23425
rect 24751 23360 24757 23424
rect 24821 23360 24837 23424
rect 24901 23360 24917 23424
rect 24981 23360 24997 23424
rect 25061 23360 25067 23424
rect 24751 23359 25067 23360
rect 34273 23424 34589 23425
rect 34273 23360 34279 23424
rect 34343 23360 34359 23424
rect 34423 23360 34439 23424
rect 34503 23360 34519 23424
rect 34583 23360 34589 23424
rect 34273 23359 34589 23360
rect 25630 22884 25636 22948
rect 25700 22946 25706 22948
rect 26417 22946 26483 22949
rect 25700 22944 26483 22946
rect 25700 22888 26422 22944
rect 26478 22888 26483 22944
rect 25700 22886 26483 22888
rect 25700 22884 25706 22886
rect 26417 22883 26483 22886
rect 10468 22880 10784 22881
rect 10468 22816 10474 22880
rect 10538 22816 10554 22880
rect 10618 22816 10634 22880
rect 10698 22816 10714 22880
rect 10778 22816 10784 22880
rect 10468 22815 10784 22816
rect 19990 22880 20306 22881
rect 19990 22816 19996 22880
rect 20060 22816 20076 22880
rect 20140 22816 20156 22880
rect 20220 22816 20236 22880
rect 20300 22816 20306 22880
rect 19990 22815 20306 22816
rect 29512 22880 29828 22881
rect 29512 22816 29518 22880
rect 29582 22816 29598 22880
rect 29662 22816 29678 22880
rect 29742 22816 29758 22880
rect 29822 22816 29828 22880
rect 29512 22815 29828 22816
rect 39034 22880 39350 22881
rect 39034 22816 39040 22880
rect 39104 22816 39120 22880
rect 39184 22816 39200 22880
rect 39264 22816 39280 22880
rect 39344 22816 39350 22880
rect 39034 22815 39350 22816
rect 0 22538 800 22568
rect 933 22538 999 22541
rect 0 22536 999 22538
rect 0 22480 938 22536
rect 994 22480 999 22536
rect 0 22478 999 22480
rect 0 22448 800 22478
rect 933 22475 999 22478
rect 39566 22448 40366 22568
rect 30230 22340 30236 22404
rect 30300 22402 30306 22404
rect 31385 22402 31451 22405
rect 30300 22400 31451 22402
rect 30300 22344 31390 22400
rect 31446 22344 31451 22400
rect 30300 22342 31451 22344
rect 30300 22340 30306 22342
rect 31385 22339 31451 22342
rect 5707 22336 6023 22337
rect 5707 22272 5713 22336
rect 5777 22272 5793 22336
rect 5857 22272 5873 22336
rect 5937 22272 5953 22336
rect 6017 22272 6023 22336
rect 5707 22271 6023 22272
rect 15229 22336 15545 22337
rect 15229 22272 15235 22336
rect 15299 22272 15315 22336
rect 15379 22272 15395 22336
rect 15459 22272 15475 22336
rect 15539 22272 15545 22336
rect 15229 22271 15545 22272
rect 24751 22336 25067 22337
rect 24751 22272 24757 22336
rect 24821 22272 24837 22336
rect 24901 22272 24917 22336
rect 24981 22272 24997 22336
rect 25061 22272 25067 22336
rect 24751 22271 25067 22272
rect 34273 22336 34589 22337
rect 34273 22272 34279 22336
rect 34343 22272 34359 22336
rect 34423 22272 34439 22336
rect 34503 22272 34519 22336
rect 34583 22272 34589 22336
rect 34273 22271 34589 22272
rect 32765 22130 32831 22133
rect 33174 22130 33180 22132
rect 32765 22128 33180 22130
rect 32765 22072 32770 22128
rect 32826 22072 33180 22128
rect 32765 22070 33180 22072
rect 32765 22067 32831 22070
rect 33174 22068 33180 22070
rect 33244 22068 33250 22132
rect 27613 21994 27679 21997
rect 27613 21992 31770 21994
rect 27613 21936 27618 21992
rect 27674 21936 31770 21992
rect 27613 21934 31770 21936
rect 27613 21931 27679 21934
rect 31710 21858 31770 21934
rect 32857 21858 32923 21861
rect 32990 21858 32996 21860
rect 31710 21856 32996 21858
rect 31710 21800 32862 21856
rect 32918 21800 32996 21856
rect 31710 21798 32996 21800
rect 32857 21795 32923 21798
rect 32990 21796 32996 21798
rect 33060 21796 33066 21860
rect 10468 21792 10784 21793
rect 10468 21728 10474 21792
rect 10538 21728 10554 21792
rect 10618 21728 10634 21792
rect 10698 21728 10714 21792
rect 10778 21728 10784 21792
rect 10468 21727 10784 21728
rect 19990 21792 20306 21793
rect 19990 21728 19996 21792
rect 20060 21728 20076 21792
rect 20140 21728 20156 21792
rect 20220 21728 20236 21792
rect 20300 21728 20306 21792
rect 19990 21727 20306 21728
rect 29512 21792 29828 21793
rect 29512 21728 29518 21792
rect 29582 21728 29598 21792
rect 29662 21728 29678 21792
rect 29742 21728 29758 21792
rect 29822 21728 29828 21792
rect 29512 21727 29828 21728
rect 39034 21792 39350 21793
rect 39034 21728 39040 21792
rect 39104 21728 39120 21792
rect 39184 21728 39200 21792
rect 39264 21728 39280 21792
rect 39344 21728 39350 21792
rect 39034 21727 39350 21728
rect 5707 21248 6023 21249
rect 5707 21184 5713 21248
rect 5777 21184 5793 21248
rect 5857 21184 5873 21248
rect 5937 21184 5953 21248
rect 6017 21184 6023 21248
rect 5707 21183 6023 21184
rect 15229 21248 15545 21249
rect 15229 21184 15235 21248
rect 15299 21184 15315 21248
rect 15379 21184 15395 21248
rect 15459 21184 15475 21248
rect 15539 21184 15545 21248
rect 15229 21183 15545 21184
rect 24751 21248 25067 21249
rect 24751 21184 24757 21248
rect 24821 21184 24837 21248
rect 24901 21184 24917 21248
rect 24981 21184 24997 21248
rect 25061 21184 25067 21248
rect 24751 21183 25067 21184
rect 34273 21248 34589 21249
rect 34273 21184 34279 21248
rect 34343 21184 34359 21248
rect 34423 21184 34439 21248
rect 34503 21184 34519 21248
rect 34583 21184 34589 21248
rect 34273 21183 34589 21184
rect 19149 21042 19215 21045
rect 22686 21042 22692 21044
rect 19149 21040 22692 21042
rect 19149 20984 19154 21040
rect 19210 20984 22692 21040
rect 19149 20982 22692 20984
rect 19149 20979 19215 20982
rect 22686 20980 22692 20982
rect 22756 20980 22762 21044
rect 12617 20906 12683 20909
rect 12750 20906 12756 20908
rect 12617 20904 12756 20906
rect 12617 20848 12622 20904
rect 12678 20848 12756 20904
rect 12617 20846 12756 20848
rect 12617 20843 12683 20846
rect 12750 20844 12756 20846
rect 12820 20844 12826 20908
rect 17902 20708 17908 20772
rect 17972 20770 17978 20772
rect 18689 20770 18755 20773
rect 17972 20768 18755 20770
rect 17972 20712 18694 20768
rect 18750 20712 18755 20768
rect 17972 20710 18755 20712
rect 17972 20708 17978 20710
rect 18689 20707 18755 20710
rect 32765 20772 32831 20773
rect 32765 20768 32812 20772
rect 32876 20770 32882 20772
rect 32765 20712 32770 20768
rect 32765 20708 32812 20712
rect 32876 20710 32922 20770
rect 32876 20708 32882 20710
rect 32765 20707 32831 20708
rect 10468 20704 10784 20705
rect 10468 20640 10474 20704
rect 10538 20640 10554 20704
rect 10618 20640 10634 20704
rect 10698 20640 10714 20704
rect 10778 20640 10784 20704
rect 10468 20639 10784 20640
rect 19990 20704 20306 20705
rect 19990 20640 19996 20704
rect 20060 20640 20076 20704
rect 20140 20640 20156 20704
rect 20220 20640 20236 20704
rect 20300 20640 20306 20704
rect 19990 20639 20306 20640
rect 29512 20704 29828 20705
rect 29512 20640 29518 20704
rect 29582 20640 29598 20704
rect 29662 20640 29678 20704
rect 29742 20640 29758 20704
rect 29822 20640 29828 20704
rect 29512 20639 29828 20640
rect 39034 20704 39350 20705
rect 39034 20640 39040 20704
rect 39104 20640 39120 20704
rect 39184 20640 39200 20704
rect 39264 20640 39280 20704
rect 39344 20640 39350 20704
rect 39034 20639 39350 20640
rect 0 20498 800 20528
rect 933 20498 999 20501
rect 0 20496 999 20498
rect 0 20440 938 20496
rect 994 20440 999 20496
rect 0 20438 999 20440
rect 0 20408 800 20438
rect 933 20435 999 20438
rect 39389 20498 39455 20501
rect 39566 20498 40366 20528
rect 39389 20496 40366 20498
rect 39389 20440 39394 20496
rect 39450 20440 40366 20496
rect 39389 20438 40366 20440
rect 39389 20435 39455 20438
rect 39566 20408 40366 20438
rect 13721 20362 13787 20365
rect 21265 20362 21331 20365
rect 13721 20360 21331 20362
rect 13721 20304 13726 20360
rect 13782 20304 21270 20360
rect 21326 20304 21331 20360
rect 13721 20302 21331 20304
rect 13721 20299 13787 20302
rect 21265 20299 21331 20302
rect 5707 20160 6023 20161
rect 5707 20096 5713 20160
rect 5777 20096 5793 20160
rect 5857 20096 5873 20160
rect 5937 20096 5953 20160
rect 6017 20096 6023 20160
rect 5707 20095 6023 20096
rect 15229 20160 15545 20161
rect 15229 20096 15235 20160
rect 15299 20096 15315 20160
rect 15379 20096 15395 20160
rect 15459 20096 15475 20160
rect 15539 20096 15545 20160
rect 15229 20095 15545 20096
rect 24751 20160 25067 20161
rect 24751 20096 24757 20160
rect 24821 20096 24837 20160
rect 24901 20096 24917 20160
rect 24981 20096 24997 20160
rect 25061 20096 25067 20160
rect 24751 20095 25067 20096
rect 34273 20160 34589 20161
rect 34273 20096 34279 20160
rect 34343 20096 34359 20160
rect 34423 20096 34439 20160
rect 34503 20096 34519 20160
rect 34583 20096 34589 20160
rect 34273 20095 34589 20096
rect 21817 20090 21883 20093
rect 23565 20090 23631 20093
rect 25773 20090 25839 20093
rect 30189 20090 30255 20093
rect 21817 20088 23631 20090
rect 21817 20032 21822 20088
rect 21878 20032 23570 20088
rect 23626 20032 23631 20088
rect 21817 20030 23631 20032
rect 21817 20027 21883 20030
rect 23565 20027 23631 20030
rect 25638 20088 30255 20090
rect 25638 20032 25778 20088
rect 25834 20032 30194 20088
rect 30250 20032 30255 20088
rect 25638 20030 30255 20032
rect 19333 19954 19399 19957
rect 21725 19954 21791 19957
rect 22185 19954 22251 19957
rect 19333 19952 19442 19954
rect 19333 19896 19338 19952
rect 19394 19896 19442 19952
rect 19333 19891 19442 19896
rect 21725 19952 22251 19954
rect 21725 19896 21730 19952
rect 21786 19896 22190 19952
rect 22246 19896 22251 19952
rect 21725 19894 22251 19896
rect 21725 19891 21791 19894
rect 22185 19891 22251 19894
rect 22829 19954 22895 19957
rect 25638 19954 25698 20030
rect 25773 20027 25839 20030
rect 30189 20027 30255 20030
rect 22829 19952 25698 19954
rect 22829 19896 22834 19952
rect 22890 19896 25698 19952
rect 22829 19894 25698 19896
rect 25865 19954 25931 19957
rect 38469 19954 38535 19957
rect 25865 19952 38535 19954
rect 25865 19896 25870 19952
rect 25926 19896 38474 19952
rect 38530 19896 38535 19952
rect 25865 19894 38535 19896
rect 22829 19891 22895 19894
rect 25865 19891 25931 19894
rect 38469 19891 38535 19894
rect 19382 19685 19442 19891
rect 19885 19818 19951 19821
rect 33685 19818 33751 19821
rect 19885 19816 33751 19818
rect 19885 19760 19890 19816
rect 19946 19760 33690 19816
rect 33746 19760 33751 19816
rect 19885 19758 33751 19760
rect 19885 19755 19951 19758
rect 33685 19755 33751 19758
rect 13629 19682 13695 19685
rect 14958 19682 14964 19684
rect 13629 19680 14964 19682
rect 13629 19624 13634 19680
rect 13690 19624 14964 19680
rect 13629 19622 14964 19624
rect 13629 19619 13695 19622
rect 14958 19620 14964 19622
rect 15028 19620 15034 19684
rect 19333 19680 19442 19685
rect 19333 19624 19338 19680
rect 19394 19624 19442 19680
rect 19333 19622 19442 19624
rect 20713 19682 20779 19685
rect 26417 19682 26483 19685
rect 20713 19680 26483 19682
rect 20713 19624 20718 19680
rect 20774 19624 26422 19680
rect 26478 19624 26483 19680
rect 20713 19622 26483 19624
rect 19333 19619 19399 19622
rect 20713 19619 20779 19622
rect 26417 19619 26483 19622
rect 10468 19616 10784 19617
rect 10468 19552 10474 19616
rect 10538 19552 10554 19616
rect 10618 19552 10634 19616
rect 10698 19552 10714 19616
rect 10778 19552 10784 19616
rect 10468 19551 10784 19552
rect 19990 19616 20306 19617
rect 19990 19552 19996 19616
rect 20060 19552 20076 19616
rect 20140 19552 20156 19616
rect 20220 19552 20236 19616
rect 20300 19552 20306 19616
rect 19990 19551 20306 19552
rect 29512 19616 29828 19617
rect 29512 19552 29518 19616
rect 29582 19552 29598 19616
rect 29662 19552 29678 19616
rect 29742 19552 29758 19616
rect 29822 19552 29828 19616
rect 29512 19551 29828 19552
rect 39034 19616 39350 19617
rect 39034 19552 39040 19616
rect 39104 19552 39120 19616
rect 39184 19552 39200 19616
rect 39264 19552 39280 19616
rect 39344 19552 39350 19616
rect 39034 19551 39350 19552
rect 13445 19546 13511 19549
rect 16021 19546 16087 19549
rect 13445 19544 16087 19546
rect 13445 19488 13450 19544
rect 13506 19488 16026 19544
rect 16082 19488 16087 19544
rect 13445 19486 16087 19488
rect 13445 19483 13511 19486
rect 16021 19483 16087 19486
rect 22093 19546 22159 19549
rect 22829 19546 22895 19549
rect 22093 19544 22895 19546
rect 22093 19488 22098 19544
rect 22154 19488 22834 19544
rect 22890 19488 22895 19544
rect 22093 19486 22895 19488
rect 22093 19483 22159 19486
rect 22829 19483 22895 19486
rect 30649 19546 30715 19549
rect 37181 19546 37247 19549
rect 30649 19544 37247 19546
rect 30649 19488 30654 19544
rect 30710 19488 37186 19544
rect 37242 19488 37247 19544
rect 30649 19486 37247 19488
rect 30649 19483 30715 19486
rect 37181 19483 37247 19486
rect 10225 19410 10291 19413
rect 14089 19410 14155 19413
rect 14273 19410 14339 19413
rect 10225 19408 14339 19410
rect 10225 19352 10230 19408
rect 10286 19352 14094 19408
rect 14150 19352 14278 19408
rect 14334 19352 14339 19408
rect 10225 19350 14339 19352
rect 10225 19347 10291 19350
rect 14089 19347 14155 19350
rect 14273 19347 14339 19350
rect 16389 19410 16455 19413
rect 24761 19410 24827 19413
rect 28349 19410 28415 19413
rect 30741 19410 30807 19413
rect 16389 19408 24827 19410
rect 16389 19352 16394 19408
rect 16450 19352 24766 19408
rect 24822 19352 24827 19408
rect 16389 19350 24827 19352
rect 16389 19347 16455 19350
rect 24761 19347 24827 19350
rect 26190 19408 30807 19410
rect 26190 19352 28354 19408
rect 28410 19352 30746 19408
rect 30802 19352 30807 19408
rect 26190 19350 30807 19352
rect 11053 19274 11119 19277
rect 13302 19274 13308 19276
rect 11053 19272 13308 19274
rect 11053 19216 11058 19272
rect 11114 19216 13308 19272
rect 11053 19214 13308 19216
rect 11053 19211 11119 19214
rect 13302 19212 13308 19214
rect 13372 19212 13378 19276
rect 14406 19212 14412 19276
rect 14476 19274 14482 19276
rect 26190 19274 26250 19350
rect 28349 19347 28415 19350
rect 30741 19347 30807 19350
rect 32622 19348 32628 19412
rect 32692 19410 32698 19412
rect 34697 19410 34763 19413
rect 32692 19408 34763 19410
rect 32692 19352 34702 19408
rect 34758 19352 34763 19408
rect 32692 19350 34763 19352
rect 32692 19348 32698 19350
rect 34697 19347 34763 19350
rect 14476 19214 26250 19274
rect 14476 19212 14482 19214
rect 5707 19072 6023 19073
rect 5707 19008 5713 19072
rect 5777 19008 5793 19072
rect 5857 19008 5873 19072
rect 5937 19008 5953 19072
rect 6017 19008 6023 19072
rect 5707 19007 6023 19008
rect 15229 19072 15545 19073
rect 15229 19008 15235 19072
rect 15299 19008 15315 19072
rect 15379 19008 15395 19072
rect 15459 19008 15475 19072
rect 15539 19008 15545 19072
rect 15229 19007 15545 19008
rect 24751 19072 25067 19073
rect 24751 19008 24757 19072
rect 24821 19008 24837 19072
rect 24901 19008 24917 19072
rect 24981 19008 24997 19072
rect 25061 19008 25067 19072
rect 24751 19007 25067 19008
rect 34273 19072 34589 19073
rect 34273 19008 34279 19072
rect 34343 19008 34359 19072
rect 34423 19008 34439 19072
rect 34503 19008 34519 19072
rect 34583 19008 34589 19072
rect 34273 19007 34589 19008
rect 15878 18804 15884 18868
rect 15948 18866 15954 18868
rect 30649 18866 30715 18869
rect 15948 18864 30715 18866
rect 15948 18808 30654 18864
rect 30710 18808 30715 18864
rect 15948 18806 30715 18808
rect 15948 18804 15954 18806
rect 30649 18803 30715 18806
rect 15653 18730 15719 18733
rect 16062 18730 16068 18732
rect 15653 18728 16068 18730
rect 15653 18672 15658 18728
rect 15714 18672 16068 18728
rect 15653 18670 16068 18672
rect 15653 18667 15719 18670
rect 16062 18668 16068 18670
rect 16132 18730 16138 18732
rect 23381 18730 23447 18733
rect 30649 18730 30715 18733
rect 16132 18728 30715 18730
rect 16132 18672 23386 18728
rect 23442 18672 30654 18728
rect 30710 18672 30715 18728
rect 16132 18670 30715 18672
rect 16132 18668 16138 18670
rect 23381 18667 23447 18670
rect 30649 18667 30715 18670
rect 25405 18596 25471 18597
rect 25405 18594 25452 18596
rect 25360 18592 25452 18594
rect 25360 18536 25410 18592
rect 25360 18534 25452 18536
rect 25405 18532 25452 18534
rect 25516 18532 25522 18596
rect 25405 18531 25471 18532
rect 10468 18528 10784 18529
rect 0 18458 800 18488
rect 10468 18464 10474 18528
rect 10538 18464 10554 18528
rect 10618 18464 10634 18528
rect 10698 18464 10714 18528
rect 10778 18464 10784 18528
rect 10468 18463 10784 18464
rect 19990 18528 20306 18529
rect 19990 18464 19996 18528
rect 20060 18464 20076 18528
rect 20140 18464 20156 18528
rect 20220 18464 20236 18528
rect 20300 18464 20306 18528
rect 19990 18463 20306 18464
rect 29512 18528 29828 18529
rect 29512 18464 29518 18528
rect 29582 18464 29598 18528
rect 29662 18464 29678 18528
rect 29742 18464 29758 18528
rect 29822 18464 29828 18528
rect 29512 18463 29828 18464
rect 39034 18528 39350 18529
rect 39034 18464 39040 18528
rect 39104 18464 39120 18528
rect 39184 18464 39200 18528
rect 39264 18464 39280 18528
rect 39344 18464 39350 18528
rect 39034 18463 39350 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 39566 18368 40366 18488
rect 6913 18322 6979 18325
rect 17401 18322 17467 18325
rect 6913 18320 17467 18322
rect 6913 18264 6918 18320
rect 6974 18264 17406 18320
rect 17462 18264 17467 18320
rect 6913 18262 17467 18264
rect 6913 18259 6979 18262
rect 17401 18259 17467 18262
rect 22318 18260 22324 18324
rect 22388 18322 22394 18324
rect 29085 18322 29151 18325
rect 22388 18320 29151 18322
rect 22388 18264 29090 18320
rect 29146 18264 29151 18320
rect 22388 18262 29151 18264
rect 22388 18260 22394 18262
rect 29085 18259 29151 18262
rect 15101 18186 15167 18189
rect 16982 18186 16988 18188
rect 15101 18184 16988 18186
rect 15101 18128 15106 18184
rect 15162 18128 16988 18184
rect 15101 18126 16988 18128
rect 15101 18123 15167 18126
rect 16982 18124 16988 18126
rect 17052 18124 17058 18188
rect 17718 18124 17724 18188
rect 17788 18186 17794 18188
rect 17861 18186 17927 18189
rect 17788 18184 17927 18186
rect 17788 18128 17866 18184
rect 17922 18128 17927 18184
rect 17788 18126 17927 18128
rect 17788 18124 17794 18126
rect 17861 18123 17927 18126
rect 26049 18186 26115 18189
rect 33726 18186 33732 18188
rect 26049 18184 33732 18186
rect 26049 18128 26054 18184
rect 26110 18128 33732 18184
rect 26049 18126 33732 18128
rect 26049 18123 26115 18126
rect 33726 18124 33732 18126
rect 33796 18124 33802 18188
rect 27061 18050 27127 18053
rect 27654 18050 27660 18052
rect 27061 18048 27660 18050
rect 27061 17992 27066 18048
rect 27122 17992 27660 18048
rect 27061 17990 27660 17992
rect 27061 17987 27127 17990
rect 27654 17988 27660 17990
rect 27724 17988 27730 18052
rect 5707 17984 6023 17985
rect 5707 17920 5713 17984
rect 5777 17920 5793 17984
rect 5857 17920 5873 17984
rect 5937 17920 5953 17984
rect 6017 17920 6023 17984
rect 5707 17919 6023 17920
rect 15229 17984 15545 17985
rect 15229 17920 15235 17984
rect 15299 17920 15315 17984
rect 15379 17920 15395 17984
rect 15459 17920 15475 17984
rect 15539 17920 15545 17984
rect 15229 17919 15545 17920
rect 24751 17984 25067 17985
rect 24751 17920 24757 17984
rect 24821 17920 24837 17984
rect 24901 17920 24917 17984
rect 24981 17920 24997 17984
rect 25061 17920 25067 17984
rect 24751 17919 25067 17920
rect 34273 17984 34589 17985
rect 34273 17920 34279 17984
rect 34343 17920 34359 17984
rect 34423 17920 34439 17984
rect 34503 17920 34519 17984
rect 34583 17920 34589 17984
rect 34273 17919 34589 17920
rect 27102 17852 27108 17916
rect 27172 17914 27178 17916
rect 27521 17914 27587 17917
rect 31661 17914 31727 17917
rect 27172 17912 31727 17914
rect 27172 17856 27526 17912
rect 27582 17856 31666 17912
rect 31722 17856 31727 17912
rect 27172 17854 31727 17856
rect 27172 17852 27178 17854
rect 27521 17851 27587 17854
rect 31661 17851 31727 17854
rect 8201 17778 8267 17781
rect 18270 17778 18276 17780
rect 8201 17776 18276 17778
rect 8201 17720 8206 17776
rect 8262 17720 18276 17776
rect 8201 17718 18276 17720
rect 8201 17715 8267 17718
rect 18270 17716 18276 17718
rect 18340 17716 18346 17780
rect 24945 17778 25011 17781
rect 25313 17778 25379 17781
rect 32489 17778 32555 17781
rect 24945 17776 32555 17778
rect 24945 17720 24950 17776
rect 25006 17720 25318 17776
rect 25374 17720 32494 17776
rect 32550 17720 32555 17776
rect 24945 17718 32555 17720
rect 24945 17715 25011 17718
rect 25313 17715 25379 17718
rect 32489 17715 32555 17718
rect 3417 17642 3483 17645
rect 24669 17642 24735 17645
rect 3417 17640 24735 17642
rect 3417 17584 3422 17640
rect 3478 17584 24674 17640
rect 24730 17584 24735 17640
rect 3417 17582 24735 17584
rect 3417 17579 3483 17582
rect 24669 17579 24735 17582
rect 25957 17642 26023 17645
rect 29361 17642 29427 17645
rect 33409 17642 33475 17645
rect 25957 17640 33475 17642
rect 25957 17584 25962 17640
rect 26018 17584 29366 17640
rect 29422 17584 33414 17640
rect 33470 17584 33475 17640
rect 25957 17582 33475 17584
rect 25957 17579 26023 17582
rect 29361 17579 29427 17582
rect 33409 17579 33475 17582
rect 10468 17440 10784 17441
rect 10468 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10784 17440
rect 10468 17375 10784 17376
rect 19990 17440 20306 17441
rect 19990 17376 19996 17440
rect 20060 17376 20076 17440
rect 20140 17376 20156 17440
rect 20220 17376 20236 17440
rect 20300 17376 20306 17440
rect 19990 17375 20306 17376
rect 29512 17440 29828 17441
rect 29512 17376 29518 17440
rect 29582 17376 29598 17440
rect 29662 17376 29678 17440
rect 29742 17376 29758 17440
rect 29822 17376 29828 17440
rect 29512 17375 29828 17376
rect 39034 17440 39350 17441
rect 39034 17376 39040 17440
rect 39104 17376 39120 17440
rect 39184 17376 39200 17440
rect 39264 17376 39280 17440
rect 39344 17376 39350 17440
rect 39034 17375 39350 17376
rect 19333 17370 19399 17373
rect 19558 17370 19564 17372
rect 19333 17368 19564 17370
rect 19333 17312 19338 17368
rect 19394 17312 19564 17368
rect 19333 17310 19564 17312
rect 19333 17307 19399 17310
rect 19558 17308 19564 17310
rect 19628 17308 19634 17372
rect 6494 17172 6500 17236
rect 6564 17234 6570 17236
rect 26601 17234 26667 17237
rect 6564 17232 26667 17234
rect 6564 17176 26606 17232
rect 26662 17176 26667 17232
rect 6564 17174 26667 17176
rect 6564 17172 6570 17174
rect 26601 17171 26667 17174
rect 29729 17234 29795 17237
rect 34145 17234 34211 17237
rect 29729 17232 34211 17234
rect 29729 17176 29734 17232
rect 29790 17176 34150 17232
rect 34206 17176 34211 17232
rect 29729 17174 34211 17176
rect 29729 17171 29795 17174
rect 34145 17171 34211 17174
rect 5165 17100 5231 17101
rect 5165 17098 5212 17100
rect 5120 17096 5212 17098
rect 5120 17040 5170 17096
rect 5120 17038 5212 17040
rect 5165 17036 5212 17038
rect 5276 17036 5282 17100
rect 5349 17098 5415 17101
rect 23657 17098 23723 17101
rect 26049 17098 26115 17101
rect 28441 17098 28507 17101
rect 5349 17096 23723 17098
rect 5349 17040 5354 17096
rect 5410 17040 23662 17096
rect 23718 17040 23723 17096
rect 5349 17038 23723 17040
rect 5165 17035 5231 17036
rect 5349 17035 5415 17038
rect 23657 17035 23723 17038
rect 24534 17096 28507 17098
rect 24534 17040 26054 17096
rect 26110 17040 28446 17096
rect 28502 17040 28507 17096
rect 24534 17038 28507 17040
rect 19517 16962 19583 16965
rect 24534 16962 24594 17038
rect 26049 17035 26115 17038
rect 28441 17035 28507 17038
rect 30097 17098 30163 17101
rect 31334 17098 31340 17100
rect 30097 17096 31340 17098
rect 30097 17040 30102 17096
rect 30158 17040 31340 17096
rect 30097 17038 31340 17040
rect 30097 17035 30163 17038
rect 31334 17036 31340 17038
rect 31404 17036 31410 17100
rect 31569 17098 31635 17101
rect 33133 17098 33199 17101
rect 31569 17096 33199 17098
rect 31569 17040 31574 17096
rect 31630 17040 33138 17096
rect 33194 17040 33199 17096
rect 31569 17038 33199 17040
rect 31569 17035 31635 17038
rect 33133 17035 33199 17038
rect 38653 17098 38719 17101
rect 39566 17098 40366 17128
rect 38653 17096 40366 17098
rect 38653 17040 38658 17096
rect 38714 17040 40366 17096
rect 38653 17038 40366 17040
rect 38653 17035 38719 17038
rect 39566 17008 40366 17038
rect 19517 16960 24594 16962
rect 19517 16904 19522 16960
rect 19578 16904 24594 16960
rect 19517 16902 24594 16904
rect 19517 16899 19583 16902
rect 5707 16896 6023 16897
rect 5707 16832 5713 16896
rect 5777 16832 5793 16896
rect 5857 16832 5873 16896
rect 5937 16832 5953 16896
rect 6017 16832 6023 16896
rect 5707 16831 6023 16832
rect 15229 16896 15545 16897
rect 15229 16832 15235 16896
rect 15299 16832 15315 16896
rect 15379 16832 15395 16896
rect 15459 16832 15475 16896
rect 15539 16832 15545 16896
rect 15229 16831 15545 16832
rect 24751 16896 25067 16897
rect 24751 16832 24757 16896
rect 24821 16832 24837 16896
rect 24901 16832 24917 16896
rect 24981 16832 24997 16896
rect 25061 16832 25067 16896
rect 24751 16831 25067 16832
rect 34273 16896 34589 16897
rect 34273 16832 34279 16896
rect 34343 16832 34359 16896
rect 34423 16832 34439 16896
rect 34503 16832 34519 16896
rect 34583 16832 34589 16896
rect 34273 16831 34589 16832
rect 18689 16826 18755 16829
rect 18689 16824 22110 16826
rect 18689 16768 18694 16824
rect 18750 16768 22110 16824
rect 18689 16766 22110 16768
rect 18689 16763 18755 16766
rect 2773 16692 2839 16693
rect 2773 16688 2820 16692
rect 2884 16690 2890 16692
rect 2773 16632 2778 16688
rect 2773 16628 2820 16632
rect 2884 16630 2930 16690
rect 2884 16628 2890 16630
rect 12198 16628 12204 16692
rect 12268 16690 12274 16692
rect 19374 16690 19380 16692
rect 12268 16630 19380 16690
rect 12268 16628 12274 16630
rect 19374 16628 19380 16630
rect 19444 16628 19450 16692
rect 22050 16690 22110 16766
rect 27061 16690 27127 16693
rect 30373 16690 30439 16693
rect 22050 16688 30439 16690
rect 22050 16632 27066 16688
rect 27122 16632 30378 16688
rect 30434 16632 30439 16688
rect 22050 16630 30439 16632
rect 2773 16627 2839 16628
rect 27061 16627 27127 16630
rect 30373 16627 30439 16630
rect 11145 16554 11211 16557
rect 26417 16554 26483 16557
rect 11145 16552 26483 16554
rect 11145 16496 11150 16552
rect 11206 16496 26422 16552
rect 26478 16496 26483 16552
rect 11145 16494 26483 16496
rect 11145 16491 11211 16494
rect 26417 16491 26483 16494
rect 28809 16554 28875 16557
rect 34881 16554 34947 16557
rect 28809 16552 34947 16554
rect 28809 16496 28814 16552
rect 28870 16496 34886 16552
rect 34942 16496 34947 16552
rect 28809 16494 34947 16496
rect 28809 16491 28875 16494
rect 34881 16491 34947 16494
rect 0 16418 800 16448
rect 933 16418 999 16421
rect 0 16416 999 16418
rect 0 16360 938 16416
rect 994 16360 999 16416
rect 0 16358 999 16360
rect 0 16328 800 16358
rect 933 16355 999 16358
rect 10468 16352 10784 16353
rect 10468 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10784 16352
rect 10468 16287 10784 16288
rect 19990 16352 20306 16353
rect 19990 16288 19996 16352
rect 20060 16288 20076 16352
rect 20140 16288 20156 16352
rect 20220 16288 20236 16352
rect 20300 16288 20306 16352
rect 19990 16287 20306 16288
rect 29512 16352 29828 16353
rect 29512 16288 29518 16352
rect 29582 16288 29598 16352
rect 29662 16288 29678 16352
rect 29742 16288 29758 16352
rect 29822 16288 29828 16352
rect 29512 16287 29828 16288
rect 39034 16352 39350 16353
rect 39034 16288 39040 16352
rect 39104 16288 39120 16352
rect 39184 16288 39200 16352
rect 39264 16288 39280 16352
rect 39344 16288 39350 16352
rect 39034 16287 39350 16288
rect 13813 16282 13879 16285
rect 13813 16280 17418 16282
rect 13813 16224 13818 16280
rect 13874 16224 17418 16280
rect 13813 16222 17418 16224
rect 13813 16219 13879 16222
rect 8661 16146 8727 16149
rect 17358 16146 17418 16222
rect 20069 16146 20135 16149
rect 8661 16144 17234 16146
rect 8661 16088 8666 16144
rect 8722 16088 17234 16144
rect 8661 16086 17234 16088
rect 17358 16144 20135 16146
rect 17358 16088 20074 16144
rect 20130 16088 20135 16144
rect 17358 16086 20135 16088
rect 8661 16083 8727 16086
rect 11053 16010 11119 16013
rect 13813 16010 13879 16013
rect 15193 16010 15259 16013
rect 4662 15950 6194 16010
rect 4521 15874 4587 15877
rect 4662 15874 4722 15950
rect 4521 15872 4722 15874
rect 4521 15816 4526 15872
rect 4582 15816 4722 15872
rect 4521 15814 4722 15816
rect 6134 15874 6194 15950
rect 11053 16008 13879 16010
rect 11053 15952 11058 16008
rect 11114 15952 13818 16008
rect 13874 15952 13879 16008
rect 11053 15950 13879 15952
rect 11053 15947 11119 15950
rect 13813 15947 13879 15950
rect 14046 16008 15259 16010
rect 14046 15952 15198 16008
rect 15254 15952 15259 16008
rect 14046 15950 15259 15952
rect 14046 15874 14106 15950
rect 15193 15947 15259 15950
rect 6134 15814 14106 15874
rect 17174 15874 17234 16086
rect 20069 16083 20135 16086
rect 20437 16146 20503 16149
rect 31477 16146 31543 16149
rect 20437 16144 31543 16146
rect 20437 16088 20442 16144
rect 20498 16088 31482 16144
rect 31538 16088 31543 16144
rect 20437 16086 31543 16088
rect 20437 16083 20503 16086
rect 31477 16083 31543 16086
rect 17309 16010 17375 16013
rect 28901 16010 28967 16013
rect 17309 16008 28967 16010
rect 17309 15952 17314 16008
rect 17370 15952 28906 16008
rect 28962 15952 28967 16008
rect 17309 15950 28967 15952
rect 17309 15947 17375 15950
rect 28901 15947 28967 15950
rect 31569 16010 31635 16013
rect 33685 16010 33751 16013
rect 34329 16010 34395 16013
rect 31569 16008 34395 16010
rect 31569 15952 31574 16008
rect 31630 15952 33690 16008
rect 33746 15952 34334 16008
rect 34390 15952 34395 16008
rect 31569 15950 34395 15952
rect 31569 15947 31635 15950
rect 33685 15947 33751 15950
rect 34329 15947 34395 15950
rect 23381 15874 23447 15877
rect 17174 15872 23447 15874
rect 17174 15816 23386 15872
rect 23442 15816 23447 15872
rect 17174 15814 23447 15816
rect 4521 15811 4587 15814
rect 23381 15811 23447 15814
rect 5707 15808 6023 15809
rect 5707 15744 5713 15808
rect 5777 15744 5793 15808
rect 5857 15744 5873 15808
rect 5937 15744 5953 15808
rect 6017 15744 6023 15808
rect 5707 15743 6023 15744
rect 15229 15808 15545 15809
rect 15229 15744 15235 15808
rect 15299 15744 15315 15808
rect 15379 15744 15395 15808
rect 15459 15744 15475 15808
rect 15539 15744 15545 15808
rect 15229 15743 15545 15744
rect 24751 15808 25067 15809
rect 24751 15744 24757 15808
rect 24821 15744 24837 15808
rect 24901 15744 24917 15808
rect 24981 15744 24997 15808
rect 25061 15744 25067 15808
rect 24751 15743 25067 15744
rect 34273 15808 34589 15809
rect 34273 15744 34279 15808
rect 34343 15744 34359 15808
rect 34423 15744 34439 15808
rect 34503 15744 34519 15808
rect 34583 15744 34589 15808
rect 34273 15743 34589 15744
rect 9121 15738 9187 15741
rect 12433 15738 12499 15741
rect 9121 15736 12499 15738
rect 9121 15680 9126 15736
rect 9182 15680 12438 15736
rect 12494 15680 12499 15736
rect 9121 15678 12499 15680
rect 9121 15675 9187 15678
rect 12433 15675 12499 15678
rect 12709 15738 12775 15741
rect 14549 15738 14615 15741
rect 12709 15736 14615 15738
rect 12709 15680 12714 15736
rect 12770 15680 14554 15736
rect 14610 15680 14615 15736
rect 12709 15678 14615 15680
rect 12709 15675 12775 15678
rect 14549 15675 14615 15678
rect 2037 15602 2103 15605
rect 24853 15602 24919 15605
rect 35433 15602 35499 15605
rect 2037 15600 24919 15602
rect 2037 15544 2042 15600
rect 2098 15544 24858 15600
rect 24914 15544 24919 15600
rect 2037 15542 24919 15544
rect 2037 15539 2103 15542
rect 24853 15539 24919 15542
rect 25086 15600 35499 15602
rect 25086 15544 35438 15600
rect 35494 15544 35499 15600
rect 25086 15542 35499 15544
rect 4337 15466 4403 15469
rect 22553 15466 22619 15469
rect 25086 15466 25146 15542
rect 35433 15539 35499 15542
rect 4337 15464 22110 15466
rect 4337 15408 4342 15464
rect 4398 15408 22110 15464
rect 4337 15406 22110 15408
rect 4337 15403 4403 15406
rect 3049 15330 3115 15333
rect 3182 15330 3188 15332
rect 3049 15328 3188 15330
rect 3049 15272 3054 15328
rect 3110 15272 3188 15328
rect 3049 15270 3188 15272
rect 3049 15267 3115 15270
rect 3182 15268 3188 15270
rect 3252 15268 3258 15332
rect 4102 15268 4108 15332
rect 4172 15330 4178 15332
rect 4797 15330 4863 15333
rect 4172 15328 4863 15330
rect 4172 15272 4802 15328
rect 4858 15272 4863 15328
rect 4172 15270 4863 15272
rect 4172 15268 4178 15270
rect 4797 15267 4863 15270
rect 6637 15330 6703 15333
rect 8293 15330 8359 15333
rect 6637 15328 8359 15330
rect 6637 15272 6642 15328
rect 6698 15272 8298 15328
rect 8354 15272 8359 15328
rect 6637 15270 8359 15272
rect 6637 15267 6703 15270
rect 8293 15267 8359 15270
rect 11329 15330 11395 15333
rect 17309 15330 17375 15333
rect 11329 15328 17375 15330
rect 11329 15272 11334 15328
rect 11390 15272 17314 15328
rect 17370 15272 17375 15328
rect 11329 15270 17375 15272
rect 22050 15330 22110 15406
rect 22553 15464 25146 15466
rect 22553 15408 22558 15464
rect 22614 15408 25146 15464
rect 22553 15406 25146 15408
rect 28901 15466 28967 15469
rect 30465 15466 30531 15469
rect 28901 15464 30531 15466
rect 28901 15408 28906 15464
rect 28962 15408 30470 15464
rect 30526 15408 30531 15464
rect 28901 15406 30531 15408
rect 22553 15403 22619 15406
rect 28901 15403 28967 15406
rect 30465 15403 30531 15406
rect 25681 15330 25747 15333
rect 29177 15330 29243 15333
rect 22050 15328 29243 15330
rect 22050 15272 25686 15328
rect 25742 15272 29182 15328
rect 29238 15272 29243 15328
rect 22050 15270 29243 15272
rect 11329 15267 11395 15270
rect 17309 15267 17375 15270
rect 25681 15267 25747 15270
rect 29177 15267 29243 15270
rect 10468 15264 10784 15265
rect 10468 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10784 15264
rect 10468 15199 10784 15200
rect 19990 15264 20306 15265
rect 19990 15200 19996 15264
rect 20060 15200 20076 15264
rect 20140 15200 20156 15264
rect 20220 15200 20236 15264
rect 20300 15200 20306 15264
rect 19990 15199 20306 15200
rect 29512 15264 29828 15265
rect 29512 15200 29518 15264
rect 29582 15200 29598 15264
rect 29662 15200 29678 15264
rect 29742 15200 29758 15264
rect 29822 15200 29828 15264
rect 29512 15199 29828 15200
rect 39034 15264 39350 15265
rect 39034 15200 39040 15264
rect 39104 15200 39120 15264
rect 39184 15200 39200 15264
rect 39264 15200 39280 15264
rect 39344 15200 39350 15264
rect 39034 15199 39350 15200
rect 2681 15194 2747 15197
rect 8477 15194 8543 15197
rect 2681 15192 8543 15194
rect 2681 15136 2686 15192
rect 2742 15136 8482 15192
rect 8538 15136 8543 15192
rect 2681 15134 8543 15136
rect 2681 15131 2747 15134
rect 8477 15131 8543 15134
rect 12065 15194 12131 15197
rect 15561 15194 15627 15197
rect 16430 15194 16436 15196
rect 12065 15192 16436 15194
rect 12065 15136 12070 15192
rect 12126 15136 15566 15192
rect 15622 15136 16436 15192
rect 12065 15134 16436 15136
rect 12065 15131 12131 15134
rect 15561 15131 15627 15134
rect 16430 15132 16436 15134
rect 16500 15132 16506 15196
rect 19374 15132 19380 15196
rect 19444 15194 19450 15196
rect 19701 15194 19767 15197
rect 19444 15192 19767 15194
rect 19444 15136 19706 15192
rect 19762 15136 19767 15192
rect 19444 15134 19767 15136
rect 19444 15132 19450 15134
rect 19701 15131 19767 15134
rect 21357 15194 21423 15197
rect 27470 15194 27476 15196
rect 21357 15192 27476 15194
rect 21357 15136 21362 15192
rect 21418 15136 27476 15192
rect 21357 15134 27476 15136
rect 21357 15131 21423 15134
rect 27470 15132 27476 15134
rect 27540 15132 27546 15196
rect 0 15058 800 15088
rect 933 15058 999 15061
rect 0 15056 999 15058
rect 0 15000 938 15056
rect 994 15000 999 15056
rect 0 14998 999 15000
rect 0 14968 800 14998
rect 933 14995 999 14998
rect 4889 15058 4955 15061
rect 11881 15058 11947 15061
rect 4889 15056 11947 15058
rect 4889 15000 4894 15056
rect 4950 15000 11886 15056
rect 11942 15000 11947 15056
rect 4889 14998 11947 15000
rect 4889 14995 4955 14998
rect 11881 14995 11947 14998
rect 12157 15058 12223 15061
rect 12934 15058 12940 15060
rect 12157 15056 12940 15058
rect 12157 15000 12162 15056
rect 12218 15000 12940 15056
rect 12157 14998 12940 15000
rect 12157 14995 12223 14998
rect 12934 14996 12940 14998
rect 13004 14996 13010 15060
rect 13261 15058 13327 15061
rect 14273 15058 14339 15061
rect 17401 15058 17467 15061
rect 13261 15056 17467 15058
rect 13261 15000 13266 15056
rect 13322 15000 14278 15056
rect 14334 15000 17406 15056
rect 17462 15000 17467 15056
rect 13261 14998 17467 15000
rect 13261 14995 13327 14998
rect 14273 14995 14339 14998
rect 17401 14995 17467 14998
rect 19558 14996 19564 15060
rect 19628 15058 19634 15060
rect 19977 15058 20043 15061
rect 19628 15056 20043 15058
rect 19628 15000 19982 15056
rect 20038 15000 20043 15056
rect 19628 14998 20043 15000
rect 19628 14996 19634 14998
rect 19977 14995 20043 14998
rect 23381 15058 23447 15061
rect 35157 15058 35223 15061
rect 23381 15056 35223 15058
rect 23381 15000 23386 15056
rect 23442 15000 35162 15056
rect 35218 15000 35223 15056
rect 23381 14998 35223 15000
rect 23381 14995 23447 14998
rect 35157 14995 35223 14998
rect 38653 15058 38719 15061
rect 39566 15058 40366 15088
rect 38653 15056 40366 15058
rect 38653 15000 38658 15056
rect 38714 15000 40366 15056
rect 38653 14998 40366 15000
rect 38653 14995 38719 14998
rect 39566 14968 40366 14998
rect 10317 14922 10383 14925
rect 17493 14922 17559 14925
rect 10317 14920 17559 14922
rect 10317 14864 10322 14920
rect 10378 14864 17498 14920
rect 17554 14864 17559 14920
rect 10317 14862 17559 14864
rect 10317 14859 10383 14862
rect 17493 14859 17559 14862
rect 19425 14922 19491 14925
rect 24117 14922 24183 14925
rect 25129 14922 25195 14925
rect 19425 14920 25195 14922
rect 19425 14864 19430 14920
rect 19486 14864 24122 14920
rect 24178 14864 25134 14920
rect 25190 14864 25195 14920
rect 19425 14862 25195 14864
rect 19425 14859 19491 14862
rect 24117 14859 24183 14862
rect 25129 14859 25195 14862
rect 16021 14786 16087 14789
rect 18505 14786 18571 14789
rect 20662 14786 20668 14788
rect 16021 14784 20668 14786
rect 16021 14728 16026 14784
rect 16082 14728 18510 14784
rect 18566 14728 20668 14784
rect 16021 14726 20668 14728
rect 16021 14723 16087 14726
rect 18505 14723 18571 14726
rect 20662 14724 20668 14726
rect 20732 14724 20738 14788
rect 5707 14720 6023 14721
rect 5707 14656 5713 14720
rect 5777 14656 5793 14720
rect 5857 14656 5873 14720
rect 5937 14656 5953 14720
rect 6017 14656 6023 14720
rect 5707 14655 6023 14656
rect 15229 14720 15545 14721
rect 15229 14656 15235 14720
rect 15299 14656 15315 14720
rect 15379 14656 15395 14720
rect 15459 14656 15475 14720
rect 15539 14656 15545 14720
rect 15229 14655 15545 14656
rect 24751 14720 25067 14721
rect 24751 14656 24757 14720
rect 24821 14656 24837 14720
rect 24901 14656 24917 14720
rect 24981 14656 24997 14720
rect 25061 14656 25067 14720
rect 24751 14655 25067 14656
rect 34273 14720 34589 14721
rect 34273 14656 34279 14720
rect 34343 14656 34359 14720
rect 34423 14656 34439 14720
rect 34503 14656 34519 14720
rect 34583 14656 34589 14720
rect 34273 14655 34589 14656
rect 10869 14650 10935 14653
rect 11789 14650 11855 14653
rect 15101 14650 15167 14653
rect 10869 14648 15167 14650
rect 10869 14592 10874 14648
rect 10930 14592 11794 14648
rect 11850 14592 15106 14648
rect 15162 14592 15167 14648
rect 10869 14590 15167 14592
rect 10869 14587 10935 14590
rect 11789 14587 11855 14590
rect 15101 14587 15167 14590
rect 4981 14514 5047 14517
rect 7097 14514 7163 14517
rect 4981 14512 7163 14514
rect 4981 14456 4986 14512
rect 5042 14456 7102 14512
rect 7158 14456 7163 14512
rect 4981 14454 7163 14456
rect 4981 14451 5047 14454
rect 7097 14451 7163 14454
rect 13813 14514 13879 14517
rect 16665 14514 16731 14517
rect 13813 14512 16731 14514
rect 13813 14456 13818 14512
rect 13874 14456 16670 14512
rect 16726 14456 16731 14512
rect 13813 14454 16731 14456
rect 13813 14451 13879 14454
rect 16665 14451 16731 14454
rect 24669 14514 24735 14517
rect 37365 14514 37431 14517
rect 24669 14512 37431 14514
rect 24669 14456 24674 14512
rect 24730 14456 37370 14512
rect 37426 14456 37431 14512
rect 24669 14454 37431 14456
rect 24669 14451 24735 14454
rect 37365 14451 37431 14454
rect 12433 14378 12499 14381
rect 13261 14378 13327 14381
rect 17861 14378 17927 14381
rect 36629 14378 36695 14381
rect 12433 14376 12634 14378
rect 12433 14320 12438 14376
rect 12494 14320 12634 14376
rect 12433 14318 12634 14320
rect 12433 14315 12499 14318
rect 12574 14242 12634 14318
rect 13261 14376 17927 14378
rect 13261 14320 13266 14376
rect 13322 14320 17866 14376
rect 17922 14320 17927 14376
rect 13261 14318 17927 14320
rect 13261 14315 13327 14318
rect 17861 14315 17927 14318
rect 18094 14376 36695 14378
rect 18094 14320 36634 14376
rect 36690 14320 36695 14376
rect 18094 14318 36695 14320
rect 13445 14242 13511 14245
rect 18094 14242 18154 14318
rect 36629 14315 36695 14318
rect 12574 14240 18154 14242
rect 12574 14184 13450 14240
rect 13506 14184 18154 14240
rect 12574 14182 18154 14184
rect 13445 14179 13511 14182
rect 10468 14176 10784 14177
rect 10468 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10784 14176
rect 10468 14111 10784 14112
rect 19990 14176 20306 14177
rect 19990 14112 19996 14176
rect 20060 14112 20076 14176
rect 20140 14112 20156 14176
rect 20220 14112 20236 14176
rect 20300 14112 20306 14176
rect 19990 14111 20306 14112
rect 29512 14176 29828 14177
rect 29512 14112 29518 14176
rect 29582 14112 29598 14176
rect 29662 14112 29678 14176
rect 29742 14112 29758 14176
rect 29822 14112 29828 14176
rect 29512 14111 29828 14112
rect 39034 14176 39350 14177
rect 39034 14112 39040 14176
rect 39104 14112 39120 14176
rect 39184 14112 39200 14176
rect 39264 14112 39280 14176
rect 39344 14112 39350 14176
rect 39034 14111 39350 14112
rect 12341 14106 12407 14109
rect 18597 14106 18663 14109
rect 12341 14104 18663 14106
rect 12341 14048 12346 14104
rect 12402 14048 18602 14104
rect 18658 14048 18663 14104
rect 12341 14046 18663 14048
rect 12341 14043 12407 14046
rect 18597 14043 18663 14046
rect 6729 13970 6795 13973
rect 8017 13970 8083 13973
rect 6729 13968 8083 13970
rect 6729 13912 6734 13968
rect 6790 13912 8022 13968
rect 8078 13912 8083 13968
rect 6729 13910 8083 13912
rect 6729 13907 6795 13910
rect 8017 13907 8083 13910
rect 8201 13970 8267 13973
rect 12566 13970 12572 13972
rect 8201 13968 12572 13970
rect 8201 13912 8206 13968
rect 8262 13912 12572 13968
rect 8201 13910 12572 13912
rect 8201 13907 8267 13910
rect 12566 13908 12572 13910
rect 12636 13908 12642 13972
rect 14089 13970 14155 13973
rect 14590 13970 14596 13972
rect 14089 13968 14596 13970
rect 14089 13912 14094 13968
rect 14150 13912 14596 13968
rect 14089 13910 14596 13912
rect 14089 13907 14155 13910
rect 14590 13908 14596 13910
rect 14660 13908 14666 13972
rect 1669 13834 1735 13837
rect 7465 13834 7531 13837
rect 26785 13834 26851 13837
rect 1669 13832 7531 13834
rect 1669 13776 1674 13832
rect 1730 13776 7470 13832
rect 7526 13776 7531 13832
rect 1669 13774 7531 13776
rect 1669 13771 1735 13774
rect 7465 13771 7531 13774
rect 9630 13832 26851 13834
rect 9630 13776 26790 13832
rect 26846 13776 26851 13832
rect 9630 13774 26851 13776
rect 6637 13698 6703 13701
rect 9630 13698 9690 13774
rect 26785 13771 26851 13774
rect 6637 13696 9690 13698
rect 6637 13640 6642 13696
rect 6698 13640 9690 13696
rect 6637 13638 9690 13640
rect 16573 13698 16639 13701
rect 16798 13698 16804 13700
rect 16573 13696 16804 13698
rect 16573 13640 16578 13696
rect 16634 13640 16804 13696
rect 16573 13638 16804 13640
rect 6637 13635 6703 13638
rect 16573 13635 16639 13638
rect 16798 13636 16804 13638
rect 16868 13636 16874 13700
rect 28993 13698 29059 13701
rect 33041 13698 33107 13701
rect 28993 13696 33107 13698
rect 28993 13640 28998 13696
rect 29054 13640 33046 13696
rect 33102 13640 33107 13696
rect 28993 13638 33107 13640
rect 28993 13635 29059 13638
rect 33041 13635 33107 13638
rect 5707 13632 6023 13633
rect 5707 13568 5713 13632
rect 5777 13568 5793 13632
rect 5857 13568 5873 13632
rect 5937 13568 5953 13632
rect 6017 13568 6023 13632
rect 5707 13567 6023 13568
rect 15229 13632 15545 13633
rect 15229 13568 15235 13632
rect 15299 13568 15315 13632
rect 15379 13568 15395 13632
rect 15459 13568 15475 13632
rect 15539 13568 15545 13632
rect 15229 13567 15545 13568
rect 24751 13632 25067 13633
rect 24751 13568 24757 13632
rect 24821 13568 24837 13632
rect 24901 13568 24917 13632
rect 24981 13568 24997 13632
rect 25061 13568 25067 13632
rect 24751 13567 25067 13568
rect 34273 13632 34589 13633
rect 34273 13568 34279 13632
rect 34343 13568 34359 13632
rect 34423 13568 34439 13632
rect 34503 13568 34519 13632
rect 34583 13568 34589 13632
rect 34273 13567 34589 13568
rect 14641 13562 14707 13565
rect 14774 13562 14780 13564
rect 14641 13560 14780 13562
rect 14641 13504 14646 13560
rect 14702 13504 14780 13560
rect 14641 13502 14780 13504
rect 14641 13499 14707 13502
rect 14774 13500 14780 13502
rect 14844 13500 14850 13564
rect 15694 13500 15700 13564
rect 15764 13562 15770 13564
rect 16757 13562 16823 13565
rect 18781 13564 18847 13565
rect 18781 13562 18828 13564
rect 15764 13560 16823 13562
rect 15764 13504 16762 13560
rect 16818 13504 16823 13560
rect 15764 13502 16823 13504
rect 18736 13560 18828 13562
rect 18736 13504 18786 13560
rect 18736 13502 18828 13504
rect 15764 13500 15770 13502
rect 16757 13499 16823 13502
rect 18781 13500 18828 13502
rect 18892 13500 18898 13564
rect 27889 13562 27955 13565
rect 28390 13562 28396 13564
rect 27889 13560 28396 13562
rect 27889 13504 27894 13560
rect 27950 13504 28396 13560
rect 27889 13502 28396 13504
rect 18781 13499 18847 13500
rect 27889 13499 27955 13502
rect 28390 13500 28396 13502
rect 28460 13500 28466 13564
rect 29085 13562 29151 13565
rect 30414 13562 30420 13564
rect 29085 13560 30420 13562
rect 29085 13504 29090 13560
rect 29146 13504 30420 13560
rect 29085 13502 30420 13504
rect 29085 13499 29151 13502
rect 30414 13500 30420 13502
rect 30484 13562 30490 13564
rect 33961 13562 34027 13565
rect 30484 13560 34027 13562
rect 30484 13504 33966 13560
rect 34022 13504 34027 13560
rect 30484 13502 34027 13504
rect 30484 13500 30490 13502
rect 33961 13499 34027 13502
rect 11605 13426 11671 13429
rect 16573 13426 16639 13429
rect 11605 13424 16639 13426
rect 11605 13368 11610 13424
rect 11666 13368 16578 13424
rect 16634 13368 16639 13424
rect 11605 13366 16639 13368
rect 11605 13363 11671 13366
rect 16573 13363 16639 13366
rect 19701 13426 19767 13429
rect 23013 13426 23079 13429
rect 19701 13424 23079 13426
rect 19701 13368 19706 13424
rect 19762 13368 23018 13424
rect 23074 13368 23079 13424
rect 19701 13366 23079 13368
rect 19701 13363 19767 13366
rect 23013 13363 23079 13366
rect 3325 13290 3391 13293
rect 13169 13290 13235 13293
rect 27838 13290 27844 13292
rect 3325 13288 12450 13290
rect 3325 13232 3330 13288
rect 3386 13232 12450 13288
rect 3325 13230 12450 13232
rect 3325 13227 3391 13230
rect 12390 13154 12450 13230
rect 13169 13288 27844 13290
rect 13169 13232 13174 13288
rect 13230 13232 27844 13288
rect 13169 13230 27844 13232
rect 13169 13227 13235 13230
rect 27838 13228 27844 13230
rect 27908 13228 27914 13292
rect 30046 13228 30052 13292
rect 30116 13290 30122 13292
rect 32857 13290 32923 13293
rect 30116 13288 32923 13290
rect 30116 13232 32862 13288
rect 32918 13232 32923 13288
rect 30116 13230 32923 13232
rect 30116 13228 30122 13230
rect 32857 13227 32923 13230
rect 16757 13154 16823 13157
rect 12390 13152 16823 13154
rect 12390 13096 16762 13152
rect 16818 13096 16823 13152
rect 12390 13094 16823 13096
rect 16757 13091 16823 13094
rect 10468 13088 10784 13089
rect 0 13018 800 13048
rect 10468 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10784 13088
rect 10468 13023 10784 13024
rect 19990 13088 20306 13089
rect 19990 13024 19996 13088
rect 20060 13024 20076 13088
rect 20140 13024 20156 13088
rect 20220 13024 20236 13088
rect 20300 13024 20306 13088
rect 19990 13023 20306 13024
rect 29512 13088 29828 13089
rect 29512 13024 29518 13088
rect 29582 13024 29598 13088
rect 29662 13024 29678 13088
rect 29742 13024 29758 13088
rect 29822 13024 29828 13088
rect 29512 13023 29828 13024
rect 39034 13088 39350 13089
rect 39034 13024 39040 13088
rect 39104 13024 39120 13088
rect 39184 13024 39200 13088
rect 39264 13024 39280 13088
rect 39344 13024 39350 13088
rect 39034 13023 39350 13024
rect 933 13018 999 13021
rect 15694 13018 15700 13020
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 12390 12958 15700 13018
rect 7281 12882 7347 12885
rect 12390 12882 12450 12958
rect 15694 12956 15700 12958
rect 15764 12956 15770 13020
rect 16389 13018 16455 13021
rect 18505 13018 18571 13021
rect 19057 13018 19123 13021
rect 16389 13016 19123 13018
rect 16389 12960 16394 13016
rect 16450 12960 18510 13016
rect 18566 12960 19062 13016
rect 19118 12960 19123 13016
rect 16389 12958 19123 12960
rect 16389 12955 16455 12958
rect 18505 12955 18571 12958
rect 19057 12955 19123 12958
rect 22001 13018 22067 13021
rect 39566 13018 40366 13048
rect 22001 13016 26986 13018
rect 22001 12960 22006 13016
rect 22062 12960 26986 13016
rect 22001 12958 26986 12960
rect 22001 12955 22067 12958
rect 7281 12880 12450 12882
rect 7281 12824 7286 12880
rect 7342 12824 12450 12880
rect 7281 12822 12450 12824
rect 13261 12882 13327 12885
rect 14457 12882 14523 12885
rect 26785 12882 26851 12885
rect 13261 12880 14523 12882
rect 13261 12824 13266 12880
rect 13322 12824 14462 12880
rect 14518 12824 14523 12880
rect 13261 12822 14523 12824
rect 7281 12819 7347 12822
rect 13261 12819 13327 12822
rect 14457 12819 14523 12822
rect 14966 12880 26851 12882
rect 14966 12824 26790 12880
rect 26846 12824 26851 12880
rect 14966 12822 26851 12824
rect 26926 12882 26986 12958
rect 39438 12958 40366 13018
rect 39438 12885 39498 12958
rect 39566 12928 40366 12958
rect 37181 12882 37247 12885
rect 26926 12880 37247 12882
rect 26926 12824 37186 12880
rect 37242 12824 37247 12880
rect 26926 12822 37247 12824
rect 7373 12746 7439 12749
rect 8017 12746 8083 12749
rect 7373 12744 8083 12746
rect 7373 12688 7378 12744
rect 7434 12688 8022 12744
rect 8078 12688 8083 12744
rect 7373 12686 8083 12688
rect 7373 12683 7439 12686
rect 8017 12683 8083 12686
rect 8886 12684 8892 12748
rect 8956 12746 8962 12748
rect 12065 12746 12131 12749
rect 12433 12746 12499 12749
rect 8956 12744 12499 12746
rect 8956 12688 12070 12744
rect 12126 12688 12438 12744
rect 12494 12688 12499 12744
rect 8956 12686 12499 12688
rect 8956 12684 8962 12686
rect 12065 12683 12131 12686
rect 12433 12683 12499 12686
rect 12709 12746 12775 12749
rect 13169 12746 13235 12749
rect 12709 12744 13235 12746
rect 12709 12688 12714 12744
rect 12770 12688 13174 12744
rect 13230 12688 13235 12744
rect 12709 12686 13235 12688
rect 12709 12683 12775 12686
rect 13169 12683 13235 12686
rect 5257 12610 5323 12613
rect 5390 12610 5396 12612
rect 5257 12608 5396 12610
rect 5257 12552 5262 12608
rect 5318 12552 5396 12608
rect 5257 12550 5396 12552
rect 5257 12547 5323 12550
rect 5390 12548 5396 12550
rect 5460 12548 5466 12612
rect 7005 12610 7071 12613
rect 7741 12610 7807 12613
rect 14966 12610 15026 12822
rect 26785 12819 26851 12822
rect 37181 12819 37247 12822
rect 39389 12880 39498 12885
rect 39389 12824 39394 12880
rect 39450 12824 39498 12880
rect 39389 12822 39498 12824
rect 39389 12819 39455 12822
rect 15101 12746 15167 12749
rect 19558 12746 19564 12748
rect 15101 12744 19564 12746
rect 15101 12688 15106 12744
rect 15162 12688 19564 12744
rect 15101 12686 19564 12688
rect 15101 12683 15167 12686
rect 19558 12684 19564 12686
rect 19628 12684 19634 12748
rect 33133 12746 33199 12749
rect 24534 12744 33199 12746
rect 24534 12688 33138 12744
rect 33194 12688 33199 12744
rect 24534 12686 33199 12688
rect 7005 12608 7114 12610
rect 7005 12552 7010 12608
rect 7066 12552 7114 12608
rect 7005 12547 7114 12552
rect 7741 12608 15026 12610
rect 7741 12552 7746 12608
rect 7802 12552 15026 12608
rect 7741 12550 15026 12552
rect 7741 12547 7807 12550
rect 15694 12548 15700 12612
rect 15764 12610 15770 12612
rect 23933 12610 23999 12613
rect 15764 12608 23999 12610
rect 15764 12552 23938 12608
rect 23994 12552 23999 12608
rect 15764 12550 23999 12552
rect 15764 12548 15770 12550
rect 23933 12547 23999 12550
rect 5707 12544 6023 12545
rect 5707 12480 5713 12544
rect 5777 12480 5793 12544
rect 5857 12480 5873 12544
rect 5937 12480 5953 12544
rect 6017 12480 6023 12544
rect 5707 12479 6023 12480
rect 7054 12474 7114 12547
rect 15229 12544 15545 12545
rect 15229 12480 15235 12544
rect 15299 12480 15315 12544
rect 15379 12480 15395 12544
rect 15459 12480 15475 12544
rect 15539 12480 15545 12544
rect 15229 12479 15545 12480
rect 13445 12474 13511 12477
rect 7054 12472 13511 12474
rect 7054 12416 13450 12472
rect 13506 12416 13511 12472
rect 7054 12414 13511 12416
rect 13445 12411 13511 12414
rect 15837 12474 15903 12477
rect 24534 12474 24594 12686
rect 33133 12683 33199 12686
rect 26969 12610 27035 12613
rect 31753 12610 31819 12613
rect 34145 12610 34211 12613
rect 26969 12608 28642 12610
rect 26969 12552 26974 12608
rect 27030 12552 28642 12608
rect 26969 12550 28642 12552
rect 26969 12547 27035 12550
rect 24751 12544 25067 12545
rect 24751 12480 24757 12544
rect 24821 12480 24837 12544
rect 24901 12480 24917 12544
rect 24981 12480 24997 12544
rect 25061 12480 25067 12544
rect 24751 12479 25067 12480
rect 15837 12472 24594 12474
rect 15837 12416 15842 12472
rect 15898 12416 24594 12472
rect 15837 12414 24594 12416
rect 28582 12474 28642 12550
rect 31753 12608 34211 12610
rect 31753 12552 31758 12608
rect 31814 12552 34150 12608
rect 34206 12552 34211 12608
rect 31753 12550 34211 12552
rect 31753 12547 31819 12550
rect 34145 12547 34211 12550
rect 34273 12544 34589 12545
rect 34273 12480 34279 12544
rect 34343 12480 34359 12544
rect 34423 12480 34439 12544
rect 34503 12480 34519 12544
rect 34583 12480 34589 12544
rect 34273 12479 34589 12480
rect 31702 12474 31708 12476
rect 28582 12414 31708 12474
rect 15837 12411 15903 12414
rect 31702 12412 31708 12414
rect 31772 12412 31778 12476
rect 33225 12474 33291 12477
rect 33777 12474 33843 12477
rect 33225 12472 33843 12474
rect 33225 12416 33230 12472
rect 33286 12416 33782 12472
rect 33838 12416 33843 12472
rect 33225 12414 33843 12416
rect 33225 12411 33291 12414
rect 33777 12411 33843 12414
rect 10225 12338 10291 12341
rect 14457 12338 14523 12341
rect 10225 12336 14523 12338
rect 10225 12280 10230 12336
rect 10286 12280 14462 12336
rect 14518 12280 14523 12336
rect 10225 12278 14523 12280
rect 10225 12275 10291 12278
rect 14457 12275 14523 12278
rect 14590 12276 14596 12340
rect 14660 12338 14666 12340
rect 15285 12338 15351 12341
rect 14660 12336 15351 12338
rect 14660 12280 15290 12336
rect 15346 12280 15351 12336
rect 14660 12278 15351 12280
rect 14660 12276 14666 12278
rect 15285 12275 15351 12278
rect 16021 12338 16087 12341
rect 16430 12338 16436 12340
rect 16021 12336 16436 12338
rect 16021 12280 16026 12336
rect 16082 12280 16436 12336
rect 16021 12278 16436 12280
rect 16021 12275 16087 12278
rect 16430 12276 16436 12278
rect 16500 12276 16506 12340
rect 17769 12338 17835 12341
rect 32029 12338 32095 12341
rect 17769 12336 32095 12338
rect 17769 12280 17774 12336
rect 17830 12280 32034 12336
rect 32090 12280 32095 12336
rect 17769 12278 32095 12280
rect 17769 12275 17835 12278
rect 32029 12275 32095 12278
rect 2773 12202 2839 12205
rect 3509 12202 3575 12205
rect 2773 12200 3575 12202
rect 2773 12144 2778 12200
rect 2834 12144 3514 12200
rect 3570 12144 3575 12200
rect 2773 12142 3575 12144
rect 2773 12139 2839 12142
rect 3509 12139 3575 12142
rect 7373 12202 7439 12205
rect 23422 12202 23428 12204
rect 7373 12200 23428 12202
rect 7373 12144 7378 12200
rect 7434 12144 23428 12200
rect 7373 12142 23428 12144
rect 7373 12139 7439 12142
rect 23422 12140 23428 12142
rect 23492 12140 23498 12204
rect 25589 12202 25655 12205
rect 31150 12202 31156 12204
rect 25589 12200 31156 12202
rect 25589 12144 25594 12200
rect 25650 12144 31156 12200
rect 25589 12142 31156 12144
rect 25589 12139 25655 12142
rect 31150 12140 31156 12142
rect 31220 12140 31226 12204
rect 9397 12068 9463 12069
rect 9397 12066 9444 12068
rect 9352 12064 9444 12066
rect 9352 12008 9402 12064
rect 9352 12006 9444 12008
rect 9397 12004 9444 12006
rect 9508 12004 9514 12068
rect 9949 12066 10015 12069
rect 10317 12066 10383 12069
rect 9949 12064 10383 12066
rect 9949 12008 9954 12064
rect 10010 12008 10322 12064
rect 10378 12008 10383 12064
rect 9949 12006 10383 12008
rect 9397 12003 9463 12004
rect 9949 12003 10015 12006
rect 10317 12003 10383 12006
rect 13854 12004 13860 12068
rect 13924 12066 13930 12068
rect 17493 12066 17559 12069
rect 13924 12064 17559 12066
rect 13924 12008 17498 12064
rect 17554 12008 17559 12064
rect 13924 12006 17559 12008
rect 13924 12004 13930 12006
rect 17493 12003 17559 12006
rect 17718 12004 17724 12068
rect 17788 12066 17794 12068
rect 17861 12066 17927 12069
rect 17788 12064 17927 12066
rect 17788 12008 17866 12064
rect 17922 12008 17927 12064
rect 17788 12006 17927 12008
rect 17788 12004 17794 12006
rect 17861 12003 17927 12006
rect 22001 12066 22067 12069
rect 22001 12064 26986 12066
rect 22001 12008 22006 12064
rect 22062 12008 26986 12064
rect 22001 12006 26986 12008
rect 22001 12003 22067 12006
rect 10468 12000 10784 12001
rect 10468 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10784 12000
rect 10468 11935 10784 11936
rect 19990 12000 20306 12001
rect 19990 11936 19996 12000
rect 20060 11936 20076 12000
rect 20140 11936 20156 12000
rect 20220 11936 20236 12000
rect 20300 11936 20306 12000
rect 19990 11935 20306 11936
rect 7005 11930 7071 11933
rect 8477 11930 8543 11933
rect 7005 11928 8543 11930
rect 7005 11872 7010 11928
rect 7066 11872 8482 11928
rect 8538 11872 8543 11928
rect 7005 11870 8543 11872
rect 7005 11867 7071 11870
rect 8477 11867 8543 11870
rect 9489 11930 9555 11933
rect 9622 11930 9628 11932
rect 9489 11928 9628 11930
rect 9489 11872 9494 11928
rect 9550 11872 9628 11928
rect 9489 11870 9628 11872
rect 9489 11867 9555 11870
rect 9622 11868 9628 11870
rect 9692 11868 9698 11932
rect 13537 11930 13603 11933
rect 17401 11930 17467 11933
rect 17677 11930 17743 11933
rect 12390 11928 17743 11930
rect 12390 11872 13542 11928
rect 13598 11872 17406 11928
rect 17462 11872 17682 11928
rect 17738 11872 17743 11928
rect 12390 11870 17743 11872
rect 8109 11794 8175 11797
rect 12390 11794 12450 11870
rect 13537 11867 13603 11870
rect 17401 11867 17467 11870
rect 17677 11867 17743 11870
rect 22185 11930 22251 11933
rect 25589 11930 25655 11933
rect 22185 11928 25655 11930
rect 22185 11872 22190 11928
rect 22246 11872 25594 11928
rect 25650 11872 25655 11928
rect 22185 11870 25655 11872
rect 22185 11867 22251 11870
rect 25589 11867 25655 11870
rect 8109 11792 12450 11794
rect 8109 11736 8114 11792
rect 8170 11736 12450 11792
rect 8109 11734 12450 11736
rect 13169 11794 13235 11797
rect 24761 11794 24827 11797
rect 25773 11796 25839 11797
rect 25773 11794 25820 11796
rect 13169 11792 24827 11794
rect 13169 11736 13174 11792
rect 13230 11736 24766 11792
rect 24822 11736 24827 11792
rect 13169 11734 24827 11736
rect 25728 11792 25820 11794
rect 25728 11736 25778 11792
rect 25728 11734 25820 11736
rect 8109 11731 8175 11734
rect 13169 11731 13235 11734
rect 24761 11731 24827 11734
rect 25773 11732 25820 11734
rect 25884 11732 25890 11796
rect 26233 11794 26299 11797
rect 26734 11794 26740 11796
rect 26233 11792 26740 11794
rect 26233 11736 26238 11792
rect 26294 11736 26740 11792
rect 26233 11734 26740 11736
rect 25773 11731 25839 11732
rect 26233 11731 26299 11734
rect 26734 11732 26740 11734
rect 26804 11732 26810 11796
rect 26926 11794 26986 12006
rect 29512 12000 29828 12001
rect 29512 11936 29518 12000
rect 29582 11936 29598 12000
rect 29662 11936 29678 12000
rect 29742 11936 29758 12000
rect 29822 11936 29828 12000
rect 29512 11935 29828 11936
rect 39034 12000 39350 12001
rect 39034 11936 39040 12000
rect 39104 11936 39120 12000
rect 39184 11936 39200 12000
rect 39264 11936 39280 12000
rect 39344 11936 39350 12000
rect 39034 11935 39350 11936
rect 30373 11930 30439 11933
rect 37089 11930 37155 11933
rect 30373 11928 37155 11930
rect 30373 11872 30378 11928
rect 30434 11872 37094 11928
rect 37150 11872 37155 11928
rect 30373 11870 37155 11872
rect 30373 11867 30439 11870
rect 37089 11867 37155 11870
rect 34973 11794 35039 11797
rect 26926 11792 35039 11794
rect 26926 11736 34978 11792
rect 35034 11736 35039 11792
rect 26926 11734 35039 11736
rect 34973 11731 35039 11734
rect 4889 11658 4955 11661
rect 5073 11658 5139 11661
rect 5809 11658 5875 11661
rect 4889 11656 5875 11658
rect 4889 11600 4894 11656
rect 4950 11600 5078 11656
rect 5134 11600 5814 11656
rect 5870 11600 5875 11656
rect 4889 11598 5875 11600
rect 4889 11595 4955 11598
rect 5073 11595 5139 11598
rect 5809 11595 5875 11598
rect 8293 11658 8359 11661
rect 17769 11658 17835 11661
rect 8293 11656 17835 11658
rect 8293 11600 8298 11656
rect 8354 11600 17774 11656
rect 17830 11600 17835 11656
rect 8293 11598 17835 11600
rect 8293 11595 8359 11598
rect 17769 11595 17835 11598
rect 23197 11658 23263 11661
rect 28206 11658 28212 11660
rect 23197 11656 28212 11658
rect 23197 11600 23202 11656
rect 23258 11600 28212 11656
rect 23197 11598 28212 11600
rect 23197 11595 23263 11598
rect 28206 11596 28212 11598
rect 28276 11658 28282 11660
rect 31201 11658 31267 11661
rect 28276 11656 31267 11658
rect 28276 11600 31206 11656
rect 31262 11600 31267 11656
rect 28276 11598 31267 11600
rect 28276 11596 28282 11598
rect 31201 11595 31267 11598
rect 8109 11522 8175 11525
rect 8293 11522 8359 11525
rect 8109 11520 8359 11522
rect 8109 11464 8114 11520
rect 8170 11464 8298 11520
rect 8354 11464 8359 11520
rect 8109 11462 8359 11464
rect 8109 11459 8175 11462
rect 8293 11459 8359 11462
rect 8477 11522 8543 11525
rect 11094 11522 11100 11524
rect 8477 11520 11100 11522
rect 8477 11464 8482 11520
rect 8538 11464 11100 11520
rect 8477 11462 11100 11464
rect 8477 11459 8543 11462
rect 11094 11460 11100 11462
rect 11164 11460 11170 11524
rect 15653 11522 15719 11525
rect 17493 11522 17559 11525
rect 15653 11520 17559 11522
rect 15653 11464 15658 11520
rect 15714 11464 17498 11520
rect 17554 11464 17559 11520
rect 15653 11462 17559 11464
rect 15653 11459 15719 11462
rect 17493 11459 17559 11462
rect 25405 11522 25471 11525
rect 28717 11522 28783 11525
rect 25405 11520 28783 11522
rect 25405 11464 25410 11520
rect 25466 11464 28722 11520
rect 28778 11464 28783 11520
rect 25405 11462 28783 11464
rect 25405 11459 25471 11462
rect 28717 11459 28783 11462
rect 33133 11522 33199 11525
rect 33317 11522 33383 11525
rect 33133 11520 33383 11522
rect 33133 11464 33138 11520
rect 33194 11464 33322 11520
rect 33378 11464 33383 11520
rect 33133 11462 33383 11464
rect 33133 11459 33199 11462
rect 33317 11459 33383 11462
rect 5707 11456 6023 11457
rect 5707 11392 5713 11456
rect 5777 11392 5793 11456
rect 5857 11392 5873 11456
rect 5937 11392 5953 11456
rect 6017 11392 6023 11456
rect 5707 11391 6023 11392
rect 15229 11456 15545 11457
rect 15229 11392 15235 11456
rect 15299 11392 15315 11456
rect 15379 11392 15395 11456
rect 15459 11392 15475 11456
rect 15539 11392 15545 11456
rect 15229 11391 15545 11392
rect 24751 11456 25067 11457
rect 24751 11392 24757 11456
rect 24821 11392 24837 11456
rect 24901 11392 24917 11456
rect 24981 11392 24997 11456
rect 25061 11392 25067 11456
rect 24751 11391 25067 11392
rect 34273 11456 34589 11457
rect 34273 11392 34279 11456
rect 34343 11392 34359 11456
rect 34423 11392 34439 11456
rect 34503 11392 34519 11456
rect 34583 11392 34589 11456
rect 34273 11391 34589 11392
rect 9806 11324 9812 11388
rect 9876 11386 9882 11388
rect 11789 11386 11855 11389
rect 15653 11386 15719 11389
rect 17861 11386 17927 11389
rect 9876 11384 15164 11386
rect 9876 11328 11794 11384
rect 11850 11328 15164 11384
rect 9876 11326 15164 11328
rect 9876 11324 9882 11326
rect 11789 11323 11855 11326
rect 1853 11250 1919 11253
rect 7598 11250 7604 11252
rect 1853 11248 7604 11250
rect 1853 11192 1858 11248
rect 1914 11192 7604 11248
rect 1853 11190 7604 11192
rect 1853 11187 1919 11190
rect 7598 11188 7604 11190
rect 7668 11188 7674 11252
rect 9857 11250 9923 11253
rect 9990 11250 9996 11252
rect 9857 11248 9996 11250
rect 9857 11192 9862 11248
rect 9918 11192 9996 11248
rect 9857 11190 9996 11192
rect 9857 11187 9923 11190
rect 9990 11188 9996 11190
rect 10060 11188 10066 11252
rect 11145 11250 11211 11253
rect 15104 11250 15164 11326
rect 15653 11384 17927 11386
rect 15653 11328 15658 11384
rect 15714 11328 17866 11384
rect 17922 11328 17927 11384
rect 15653 11326 17927 11328
rect 15653 11323 15719 11326
rect 17861 11323 17927 11326
rect 21817 11386 21883 11389
rect 22461 11386 22527 11389
rect 21817 11384 22527 11386
rect 21817 11328 21822 11384
rect 21878 11328 22466 11384
rect 22522 11328 22527 11384
rect 21817 11326 22527 11328
rect 21817 11323 21883 11326
rect 22461 11323 22527 11326
rect 25313 11386 25379 11389
rect 26141 11386 26207 11389
rect 27889 11386 27955 11389
rect 25313 11384 27955 11386
rect 25313 11328 25318 11384
rect 25374 11328 26146 11384
rect 26202 11328 27894 11384
rect 27950 11328 27955 11384
rect 25313 11326 27955 11328
rect 25313 11323 25379 11326
rect 26141 11323 26207 11326
rect 27889 11323 27955 11326
rect 23013 11250 23079 11253
rect 27521 11250 27587 11253
rect 11145 11248 15026 11250
rect 11145 11192 11150 11248
rect 11206 11192 15026 11248
rect 11145 11190 15026 11192
rect 15104 11248 23079 11250
rect 15104 11192 23018 11248
rect 23074 11192 23079 11248
rect 15104 11190 23079 11192
rect 11145 11187 11211 11190
rect 10225 11116 10291 11117
rect 10174 11114 10180 11116
rect 10134 11054 10180 11114
rect 10244 11112 10291 11116
rect 10286 11056 10291 11112
rect 10174 11052 10180 11054
rect 10244 11052 10291 11056
rect 10225 11051 10291 11052
rect 11838 11054 12266 11114
rect 0 10978 800 11008
rect 933 10978 999 10981
rect 0 10976 999 10978
rect 0 10920 938 10976
rect 994 10920 999 10976
rect 0 10918 999 10920
rect 0 10888 800 10918
rect 933 10915 999 10918
rect 10468 10912 10784 10913
rect 10468 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10784 10912
rect 10468 10847 10784 10848
rect 11838 10842 11898 11054
rect 12065 10980 12131 10981
rect 12014 10978 12020 10980
rect 11974 10918 12020 10978
rect 12084 10976 12131 10980
rect 12126 10920 12131 10976
rect 12014 10916 12020 10918
rect 12084 10916 12131 10920
rect 12206 10978 12266 11054
rect 14966 10978 15026 11190
rect 23013 11187 23079 11190
rect 23430 11248 27587 11250
rect 23430 11192 27526 11248
rect 27582 11192 27587 11248
rect 23430 11190 27587 11192
rect 15377 11114 15443 11117
rect 16062 11114 16068 11116
rect 15377 11112 16068 11114
rect 15377 11056 15382 11112
rect 15438 11056 16068 11112
rect 15377 11054 16068 11056
rect 15377 11051 15443 11054
rect 16062 11052 16068 11054
rect 16132 11052 16138 11116
rect 16573 11114 16639 11117
rect 16941 11116 17007 11117
rect 16798 11114 16804 11116
rect 16573 11112 16804 11114
rect 16573 11056 16578 11112
rect 16634 11056 16804 11112
rect 16573 11054 16804 11056
rect 16573 11051 16639 11054
rect 16798 11052 16804 11054
rect 16868 11052 16874 11116
rect 16941 11112 16988 11116
rect 17052 11114 17058 11116
rect 22921 11114 22987 11117
rect 23430 11114 23490 11190
rect 27521 11187 27587 11190
rect 16941 11056 16946 11112
rect 16941 11052 16988 11056
rect 17052 11054 17098 11114
rect 22921 11112 23490 11114
rect 22921 11056 22926 11112
rect 22982 11056 23490 11112
rect 22921 11054 23490 11056
rect 23565 11114 23631 11117
rect 25313 11114 25379 11117
rect 23565 11112 25379 11114
rect 23565 11056 23570 11112
rect 23626 11056 25318 11112
rect 25374 11056 25379 11112
rect 23565 11054 25379 11056
rect 17052 11052 17058 11054
rect 16941 11051 17007 11052
rect 22921 11051 22987 11054
rect 23565 11051 23631 11054
rect 25313 11051 25379 11054
rect 25589 11114 25655 11117
rect 27981 11114 28047 11117
rect 31201 11116 31267 11117
rect 25589 11112 28047 11114
rect 25589 11056 25594 11112
rect 25650 11056 27986 11112
rect 28042 11056 28047 11112
rect 25589 11054 28047 11056
rect 25589 11051 25655 11054
rect 27981 11051 28047 11054
rect 31150 11052 31156 11116
rect 31220 11114 31267 11116
rect 31220 11112 31312 11114
rect 31262 11056 31312 11112
rect 31220 11054 31312 11056
rect 33961 11112 34027 11117
rect 33961 11056 33966 11112
rect 34022 11056 34027 11112
rect 31220 11052 31267 11054
rect 31201 11051 31267 11052
rect 33961 11051 34027 11056
rect 39389 11114 39455 11117
rect 39389 11112 39498 11114
rect 39389 11056 39394 11112
rect 39450 11056 39498 11112
rect 39389 11051 39498 11056
rect 16205 10978 16271 10981
rect 18597 10978 18663 10981
rect 12206 10918 14842 10978
rect 14966 10976 16271 10978
rect 14966 10920 16210 10976
rect 16266 10920 16271 10976
rect 14966 10918 16271 10920
rect 12065 10915 12131 10916
rect 10918 10782 11898 10842
rect 5717 10706 5783 10709
rect 7373 10706 7439 10709
rect 5717 10704 7439 10706
rect 5717 10648 5722 10704
rect 5778 10648 7378 10704
rect 7434 10648 7439 10704
rect 5717 10646 7439 10648
rect 5717 10643 5783 10646
rect 7373 10643 7439 10646
rect 8201 10706 8267 10709
rect 10918 10706 10978 10782
rect 12934 10780 12940 10844
rect 13004 10842 13010 10844
rect 13445 10842 13511 10845
rect 14457 10844 14523 10845
rect 13004 10840 13511 10842
rect 13004 10784 13450 10840
rect 13506 10784 13511 10840
rect 13004 10782 13511 10784
rect 13004 10780 13010 10782
rect 13445 10779 13511 10782
rect 14406 10780 14412 10844
rect 14476 10842 14523 10844
rect 14782 10842 14842 10918
rect 16205 10915 16271 10918
rect 17358 10976 18663 10978
rect 17358 10920 18602 10976
rect 18658 10920 18663 10976
rect 17358 10918 18663 10920
rect 15694 10842 15700 10844
rect 14476 10840 14568 10842
rect 14518 10784 14568 10840
rect 14476 10782 14568 10784
rect 14782 10782 15700 10842
rect 14476 10780 14523 10782
rect 15694 10780 15700 10782
rect 15764 10780 15770 10844
rect 16021 10842 16087 10845
rect 17358 10842 17418 10918
rect 18597 10915 18663 10918
rect 25446 10916 25452 10980
rect 25516 10978 25522 10980
rect 25681 10978 25747 10981
rect 29310 10978 29316 10980
rect 25516 10976 25747 10978
rect 25516 10920 25686 10976
rect 25742 10920 25747 10976
rect 25516 10918 25747 10920
rect 25516 10916 25522 10918
rect 25681 10915 25747 10918
rect 26788 10918 29316 10978
rect 19990 10912 20306 10913
rect 19990 10848 19996 10912
rect 20060 10848 20076 10912
rect 20140 10848 20156 10912
rect 20220 10848 20236 10912
rect 20300 10848 20306 10912
rect 19990 10847 20306 10848
rect 26788 10842 26848 10918
rect 29310 10916 29316 10918
rect 29380 10916 29386 10980
rect 30281 10978 30347 10981
rect 33964 10978 34024 11051
rect 30281 10976 34024 10978
rect 30281 10920 30286 10976
rect 30342 10920 34024 10976
rect 30281 10918 34024 10920
rect 39438 10978 39498 11051
rect 39566 10978 40366 11008
rect 39438 10918 40366 10978
rect 30281 10915 30347 10918
rect 29512 10912 29828 10913
rect 29512 10848 29518 10912
rect 29582 10848 29598 10912
rect 29662 10848 29678 10912
rect 29742 10848 29758 10912
rect 29822 10848 29828 10912
rect 29512 10847 29828 10848
rect 39034 10912 39350 10913
rect 39034 10848 39040 10912
rect 39104 10848 39120 10912
rect 39184 10848 39200 10912
rect 39264 10848 39280 10912
rect 39344 10848 39350 10912
rect 39566 10888 40366 10918
rect 39034 10847 39350 10848
rect 27521 10844 27587 10845
rect 27470 10842 27476 10844
rect 16021 10840 17418 10842
rect 16021 10784 16026 10840
rect 16082 10784 17418 10840
rect 16021 10782 17418 10784
rect 24166 10782 26848 10842
rect 27430 10782 27476 10842
rect 27540 10840 27587 10844
rect 27582 10784 27587 10840
rect 14457 10779 14523 10780
rect 16021 10779 16087 10782
rect 8201 10704 10978 10706
rect 8201 10648 8206 10704
rect 8262 10648 10978 10704
rect 8201 10646 10978 10648
rect 11145 10706 11211 10709
rect 24166 10706 24226 10782
rect 27470 10780 27476 10782
rect 27540 10780 27587 10784
rect 27521 10779 27587 10780
rect 30741 10842 30807 10845
rect 35525 10842 35591 10845
rect 30741 10840 35591 10842
rect 30741 10784 30746 10840
rect 30802 10784 35530 10840
rect 35586 10784 35591 10840
rect 30741 10782 35591 10784
rect 30741 10779 30807 10782
rect 35525 10779 35591 10782
rect 11145 10704 24226 10706
rect 11145 10648 11150 10704
rect 11206 10648 24226 10704
rect 11145 10646 24226 10648
rect 24761 10706 24827 10709
rect 37641 10706 37707 10709
rect 24761 10704 37707 10706
rect 24761 10648 24766 10704
rect 24822 10648 37646 10704
rect 37702 10648 37707 10704
rect 24761 10646 37707 10648
rect 8201 10643 8267 10646
rect 11145 10643 11211 10646
rect 24761 10643 24827 10646
rect 37641 10643 37707 10646
rect 5441 10570 5507 10573
rect 16205 10570 16271 10573
rect 25405 10570 25471 10573
rect 5441 10568 15716 10570
rect 5441 10512 5446 10568
rect 5502 10512 15716 10568
rect 5441 10510 15716 10512
rect 5441 10507 5507 10510
rect 15656 10437 15716 10510
rect 16205 10568 25471 10570
rect 16205 10512 16210 10568
rect 16266 10512 25410 10568
rect 25466 10512 25471 10568
rect 16205 10510 25471 10512
rect 16205 10507 16271 10510
rect 25405 10507 25471 10510
rect 25589 10570 25655 10573
rect 29085 10570 29151 10573
rect 25589 10568 29151 10570
rect 25589 10512 25594 10568
rect 25650 10512 29090 10568
rect 29146 10512 29151 10568
rect 25589 10510 29151 10512
rect 25589 10507 25655 10510
rect 29085 10507 29151 10510
rect 29310 10508 29316 10572
rect 29380 10570 29386 10572
rect 29821 10570 29887 10573
rect 29380 10568 29887 10570
rect 29380 10512 29826 10568
rect 29882 10512 29887 10568
rect 29380 10510 29887 10512
rect 29380 10508 29386 10510
rect 29821 10507 29887 10510
rect 15653 10434 15719 10437
rect 22645 10434 22711 10437
rect 15653 10432 22711 10434
rect 15653 10376 15658 10432
rect 15714 10376 22650 10432
rect 22706 10376 22711 10432
rect 15653 10374 22711 10376
rect 15653 10371 15719 10374
rect 22645 10371 22711 10374
rect 25313 10434 25379 10437
rect 25589 10434 25655 10437
rect 25313 10432 25655 10434
rect 25313 10376 25318 10432
rect 25374 10376 25594 10432
rect 25650 10376 25655 10432
rect 25313 10374 25655 10376
rect 25313 10371 25379 10374
rect 25589 10371 25655 10374
rect 25865 10434 25931 10437
rect 26785 10434 26851 10437
rect 25865 10432 26851 10434
rect 25865 10376 25870 10432
rect 25926 10376 26790 10432
rect 26846 10376 26851 10432
rect 25865 10374 26851 10376
rect 25865 10371 25931 10374
rect 26785 10371 26851 10374
rect 27429 10434 27495 10437
rect 33961 10434 34027 10437
rect 27429 10432 34027 10434
rect 27429 10376 27434 10432
rect 27490 10376 33966 10432
rect 34022 10376 34027 10432
rect 27429 10374 34027 10376
rect 27429 10371 27495 10374
rect 33961 10371 34027 10374
rect 5707 10368 6023 10369
rect 5707 10304 5713 10368
rect 5777 10304 5793 10368
rect 5857 10304 5873 10368
rect 5937 10304 5953 10368
rect 6017 10304 6023 10368
rect 5707 10303 6023 10304
rect 15229 10368 15545 10369
rect 15229 10304 15235 10368
rect 15299 10304 15315 10368
rect 15379 10304 15395 10368
rect 15459 10304 15475 10368
rect 15539 10304 15545 10368
rect 15229 10303 15545 10304
rect 24751 10368 25067 10369
rect 24751 10304 24757 10368
rect 24821 10304 24837 10368
rect 24901 10304 24917 10368
rect 24981 10304 24997 10368
rect 25061 10304 25067 10368
rect 24751 10303 25067 10304
rect 34273 10368 34589 10369
rect 34273 10304 34279 10368
rect 34343 10304 34359 10368
rect 34423 10304 34439 10368
rect 34503 10304 34519 10368
rect 34583 10304 34589 10368
rect 34273 10303 34589 10304
rect 11789 10298 11855 10301
rect 12893 10298 12959 10301
rect 11789 10296 12959 10298
rect 11789 10240 11794 10296
rect 11850 10240 12898 10296
rect 12954 10240 12959 10296
rect 11789 10238 12959 10240
rect 11789 10235 11855 10238
rect 12893 10235 12959 10238
rect 15837 10298 15903 10301
rect 25129 10298 25195 10301
rect 30741 10298 30807 10301
rect 15837 10296 22110 10298
rect 15837 10240 15842 10296
rect 15898 10240 22110 10296
rect 15837 10238 22110 10240
rect 15837 10235 15903 10238
rect 9765 10162 9831 10165
rect 20713 10162 20779 10165
rect 9765 10160 20779 10162
rect 9765 10104 9770 10160
rect 9826 10104 20718 10160
rect 20774 10104 20779 10160
rect 9765 10102 20779 10104
rect 22050 10162 22110 10238
rect 25129 10296 30807 10298
rect 25129 10240 25134 10296
rect 25190 10240 30746 10296
rect 30802 10240 30807 10296
rect 25129 10238 30807 10240
rect 25129 10235 25195 10238
rect 30741 10235 30807 10238
rect 32581 10298 32647 10301
rect 33225 10298 33291 10301
rect 34053 10298 34119 10301
rect 32581 10296 34119 10298
rect 32581 10240 32586 10296
rect 32642 10240 33230 10296
rect 33286 10240 34058 10296
rect 34114 10240 34119 10296
rect 32581 10238 34119 10240
rect 32581 10235 32647 10238
rect 33225 10235 33291 10238
rect 34053 10235 34119 10238
rect 27429 10162 27495 10165
rect 22050 10160 27495 10162
rect 22050 10104 27434 10160
rect 27490 10104 27495 10160
rect 22050 10102 27495 10104
rect 9765 10099 9831 10102
rect 20713 10099 20779 10102
rect 27429 10099 27495 10102
rect 28942 10100 28948 10164
rect 29012 10162 29018 10164
rect 38193 10162 38259 10165
rect 29012 10160 38259 10162
rect 29012 10104 38198 10160
rect 38254 10104 38259 10160
rect 29012 10102 38259 10104
rect 29012 10100 29018 10102
rect 38193 10099 38259 10102
rect 2221 10026 2287 10029
rect 12525 10026 12591 10029
rect 15837 10026 15903 10029
rect 36169 10026 36235 10029
rect 2221 10024 12450 10026
rect 2221 9968 2226 10024
rect 2282 9968 12450 10024
rect 2221 9966 12450 9968
rect 2221 9963 2287 9966
rect 9765 9892 9831 9893
rect 12065 9892 12131 9893
rect 9765 9890 9812 9892
rect 9720 9888 9812 9890
rect 9720 9832 9770 9888
rect 9720 9830 9812 9832
rect 9765 9828 9812 9830
rect 9876 9828 9882 9892
rect 12014 9890 12020 9892
rect 11974 9830 12020 9890
rect 12084 9888 12131 9892
rect 12126 9832 12131 9888
rect 12014 9828 12020 9830
rect 12084 9828 12131 9832
rect 12390 9890 12450 9966
rect 12525 10024 15903 10026
rect 12525 9968 12530 10024
rect 12586 9968 15842 10024
rect 15898 9968 15903 10024
rect 12525 9966 15903 9968
rect 12525 9963 12591 9966
rect 15837 9963 15903 9966
rect 17358 9966 20546 10026
rect 17217 9890 17283 9893
rect 12390 9888 17283 9890
rect 12390 9832 17222 9888
rect 17278 9832 17283 9888
rect 12390 9830 17283 9832
rect 9765 9827 9831 9828
rect 12065 9827 12131 9828
rect 17217 9827 17283 9830
rect 10468 9824 10784 9825
rect 10468 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10784 9824
rect 10468 9759 10784 9760
rect 2589 9756 2655 9757
rect 2589 9752 2636 9756
rect 2700 9754 2706 9756
rect 6361 9754 6427 9757
rect 8293 9754 8359 9757
rect 9121 9754 9187 9757
rect 2589 9696 2594 9752
rect 2589 9692 2636 9696
rect 2700 9694 2746 9754
rect 6361 9752 9187 9754
rect 6361 9696 6366 9752
rect 6422 9696 8298 9752
rect 8354 9696 9126 9752
rect 9182 9696 9187 9752
rect 6361 9694 9187 9696
rect 2700 9692 2706 9694
rect 2589 9691 2655 9692
rect 6361 9691 6427 9694
rect 8293 9691 8359 9694
rect 9121 9691 9187 9694
rect 9857 9754 9923 9757
rect 9990 9754 9996 9756
rect 9857 9752 9996 9754
rect 9857 9696 9862 9752
rect 9918 9696 9996 9752
rect 9857 9694 9996 9696
rect 9857 9691 9923 9694
rect 9990 9692 9996 9694
rect 10060 9692 10066 9756
rect 11053 9754 11119 9757
rect 11789 9754 11855 9757
rect 17358 9754 17418 9966
rect 20486 9890 20546 9966
rect 22050 10024 36235 10026
rect 22050 9968 36174 10024
rect 36230 9968 36235 10024
rect 22050 9966 36235 9968
rect 22050 9890 22110 9966
rect 36169 9963 36235 9966
rect 20486 9830 22110 9890
rect 22277 9890 22343 9893
rect 25037 9890 25103 9893
rect 22277 9888 25103 9890
rect 22277 9832 22282 9888
rect 22338 9832 25042 9888
rect 25098 9832 25103 9888
rect 22277 9830 25103 9832
rect 22277 9827 22343 9830
rect 25037 9827 25103 9830
rect 25405 9890 25471 9893
rect 29126 9890 29132 9892
rect 25405 9888 29132 9890
rect 25405 9832 25410 9888
rect 25466 9832 29132 9888
rect 25405 9830 29132 9832
rect 25405 9827 25471 9830
rect 29126 9828 29132 9830
rect 29196 9828 29202 9892
rect 32857 9890 32923 9893
rect 35709 9890 35775 9893
rect 32857 9888 35775 9890
rect 32857 9832 32862 9888
rect 32918 9832 35714 9888
rect 35770 9832 35775 9888
rect 32857 9830 35775 9832
rect 32857 9827 32923 9830
rect 35709 9827 35775 9830
rect 19990 9824 20306 9825
rect 19990 9760 19996 9824
rect 20060 9760 20076 9824
rect 20140 9760 20156 9824
rect 20220 9760 20236 9824
rect 20300 9760 20306 9824
rect 19990 9759 20306 9760
rect 29512 9824 29828 9825
rect 29512 9760 29518 9824
rect 29582 9760 29598 9824
rect 29662 9760 29678 9824
rect 29742 9760 29758 9824
rect 29822 9760 29828 9824
rect 29512 9759 29828 9760
rect 39034 9824 39350 9825
rect 39034 9760 39040 9824
rect 39104 9760 39120 9824
rect 39184 9760 39200 9824
rect 39264 9760 39280 9824
rect 39344 9760 39350 9824
rect 39034 9759 39350 9760
rect 11053 9752 11855 9754
rect 11053 9696 11058 9752
rect 11114 9696 11794 9752
rect 11850 9696 11855 9752
rect 11053 9694 11855 9696
rect 11053 9691 11119 9694
rect 11789 9691 11855 9694
rect 12390 9694 17418 9754
rect 18689 9754 18755 9757
rect 21725 9754 21791 9757
rect 25129 9754 25195 9757
rect 18689 9752 19810 9754
rect 18689 9696 18694 9752
rect 18750 9696 19810 9752
rect 18689 9694 19810 9696
rect 10317 9618 10383 9621
rect 11881 9618 11947 9621
rect 10317 9616 11947 9618
rect 10317 9560 10322 9616
rect 10378 9560 11886 9616
rect 11942 9560 11947 9616
rect 10317 9558 11947 9560
rect 10317 9555 10383 9558
rect 11881 9555 11947 9558
rect 1761 9482 1827 9485
rect 9765 9482 9831 9485
rect 1761 9480 9831 9482
rect 1761 9424 1766 9480
rect 1822 9424 9770 9480
rect 9826 9424 9831 9480
rect 1761 9422 9831 9424
rect 1761 9419 1827 9422
rect 9765 9419 9831 9422
rect 11789 9482 11855 9485
rect 12390 9482 12450 9694
rect 18689 9691 18755 9694
rect 12525 9618 12591 9621
rect 12750 9618 12756 9620
rect 12525 9616 12756 9618
rect 12525 9560 12530 9616
rect 12586 9560 12756 9616
rect 12525 9558 12756 9560
rect 12525 9555 12591 9558
rect 12750 9556 12756 9558
rect 12820 9556 12826 9620
rect 13118 9556 13124 9620
rect 13188 9618 13194 9620
rect 13188 9584 15072 9618
rect 13188 9558 15348 9584
rect 13188 9556 13194 9558
rect 11789 9480 12450 9482
rect 11789 9424 11794 9480
rect 11850 9424 12450 9480
rect 11789 9422 12450 9424
rect 11789 9419 11855 9422
rect 10409 9346 10475 9349
rect 13126 9346 13186 9556
rect 15012 9524 15348 9558
rect 15694 9556 15700 9620
rect 15764 9618 15770 9620
rect 16021 9618 16087 9621
rect 15764 9616 16087 9618
rect 15764 9560 16026 9616
rect 16082 9560 16087 9616
rect 15764 9558 16087 9560
rect 15764 9556 15770 9558
rect 16021 9555 16087 9558
rect 16481 9618 16547 9621
rect 19517 9618 19583 9621
rect 16481 9616 19583 9618
rect 16481 9560 16486 9616
rect 16542 9560 19522 9616
rect 19578 9560 19583 9616
rect 16481 9558 19583 9560
rect 19750 9618 19810 9694
rect 21725 9752 25195 9754
rect 21725 9696 21730 9752
rect 21786 9696 25134 9752
rect 25190 9696 25195 9752
rect 21725 9694 25195 9696
rect 21725 9691 21791 9694
rect 25129 9691 25195 9694
rect 26918 9692 26924 9756
rect 26988 9754 26994 9756
rect 27153 9754 27219 9757
rect 27889 9756 27955 9757
rect 26988 9752 27219 9754
rect 26988 9696 27158 9752
rect 27214 9696 27219 9752
rect 26988 9694 27219 9696
rect 26988 9692 26994 9694
rect 27153 9691 27219 9694
rect 27838 9692 27844 9756
rect 27908 9754 27955 9756
rect 28257 9754 28323 9757
rect 30189 9756 30255 9757
rect 31385 9756 31451 9757
rect 30189 9754 30236 9756
rect 27908 9752 28000 9754
rect 27950 9696 28000 9752
rect 27908 9694 28000 9696
rect 28257 9752 29424 9754
rect 28257 9696 28262 9752
rect 28318 9696 29424 9752
rect 28257 9694 29424 9696
rect 30144 9752 30236 9754
rect 30144 9696 30194 9752
rect 30144 9694 30236 9696
rect 27908 9692 27955 9694
rect 27889 9691 27955 9692
rect 28257 9691 28323 9694
rect 19977 9618 20043 9621
rect 22277 9618 22343 9621
rect 22737 9620 22803 9621
rect 22686 9618 22692 9620
rect 19750 9616 22343 9618
rect 19750 9560 19982 9616
rect 20038 9560 22282 9616
rect 22338 9560 22343 9616
rect 19750 9558 22343 9560
rect 22646 9558 22692 9618
rect 22756 9616 22803 9620
rect 22798 9560 22803 9616
rect 16481 9555 16547 9558
rect 19517 9555 19583 9558
rect 19977 9555 20043 9558
rect 22277 9555 22343 9558
rect 22686 9556 22692 9558
rect 22756 9556 22803 9560
rect 22737 9555 22803 9556
rect 24485 9618 24551 9621
rect 27705 9618 27771 9621
rect 24485 9616 27771 9618
rect 24485 9560 24490 9616
rect 24546 9560 27710 9616
rect 27766 9560 27771 9616
rect 24485 9558 27771 9560
rect 27892 9618 27952 9691
rect 28574 9618 28580 9620
rect 27892 9558 28580 9618
rect 24485 9555 24551 9558
rect 27705 9555 27771 9558
rect 28574 9556 28580 9558
rect 28644 9556 28650 9620
rect 28717 9618 28783 9621
rect 28993 9618 29059 9621
rect 28717 9616 29059 9618
rect 28717 9560 28722 9616
rect 28778 9560 28998 9616
rect 29054 9560 29059 9616
rect 28717 9558 29059 9560
rect 29364 9618 29424 9694
rect 30189 9692 30236 9694
rect 30300 9692 30306 9756
rect 31334 9754 31340 9756
rect 31258 9694 31340 9754
rect 31404 9754 31451 9756
rect 35249 9754 35315 9757
rect 31404 9752 35315 9754
rect 31446 9696 35254 9752
rect 35310 9696 35315 9752
rect 31334 9692 31340 9694
rect 31404 9694 35315 9696
rect 31404 9692 31451 9694
rect 30189 9691 30255 9692
rect 31385 9691 31451 9692
rect 35249 9691 35315 9694
rect 30833 9618 30899 9621
rect 29364 9616 30899 9618
rect 29364 9560 30838 9616
rect 30894 9560 30899 9616
rect 29364 9558 30899 9560
rect 28717 9555 28783 9558
rect 28993 9555 29059 9558
rect 30833 9555 30899 9558
rect 31886 9556 31892 9620
rect 31956 9618 31962 9620
rect 34053 9618 34119 9621
rect 31956 9616 34119 9618
rect 31956 9560 34058 9616
rect 34114 9560 34119 9616
rect 31956 9558 34119 9560
rect 31956 9556 31962 9558
rect 34053 9555 34119 9558
rect 34513 9618 34579 9621
rect 36537 9618 36603 9621
rect 34513 9616 36603 9618
rect 34513 9560 34518 9616
rect 34574 9560 36542 9616
rect 36598 9560 36603 9616
rect 34513 9558 36603 9560
rect 34513 9555 34579 9558
rect 36537 9555 36603 9558
rect 39389 9618 39455 9621
rect 39566 9618 40366 9648
rect 39389 9616 40366 9618
rect 39389 9560 39394 9616
rect 39450 9560 40366 9616
rect 39389 9558 40366 9560
rect 39389 9555 39455 9558
rect 39566 9528 40366 9558
rect 13486 9420 13492 9484
rect 13556 9482 13562 9484
rect 14365 9482 14431 9485
rect 13556 9480 14431 9482
rect 13556 9424 14370 9480
rect 14426 9424 14431 9480
rect 13556 9422 14431 9424
rect 15288 9482 15348 9524
rect 17769 9482 17835 9485
rect 27838 9482 27844 9484
rect 15288 9422 16682 9482
rect 13556 9420 13562 9422
rect 14365 9419 14431 9422
rect 10409 9344 13186 9346
rect 10409 9288 10414 9344
rect 10470 9288 13186 9344
rect 10409 9286 13186 9288
rect 13905 9346 13971 9349
rect 14038 9346 14044 9348
rect 13905 9344 14044 9346
rect 13905 9288 13910 9344
rect 13966 9288 14044 9344
rect 13905 9286 14044 9288
rect 10409 9283 10475 9286
rect 13905 9283 13971 9286
rect 14038 9284 14044 9286
rect 14108 9284 14114 9348
rect 16622 9346 16682 9422
rect 17769 9480 27844 9482
rect 17769 9424 17774 9480
rect 17830 9424 27844 9480
rect 17769 9422 27844 9424
rect 17769 9419 17835 9422
rect 27838 9420 27844 9422
rect 27908 9420 27914 9484
rect 28022 9420 28028 9484
rect 28092 9482 28098 9484
rect 28993 9482 29059 9485
rect 28092 9480 29059 9482
rect 28092 9424 28998 9480
rect 29054 9424 29059 9480
rect 28092 9422 29059 9424
rect 28092 9420 28098 9422
rect 28993 9419 29059 9422
rect 19057 9346 19123 9349
rect 21081 9346 21147 9349
rect 16622 9344 21147 9346
rect 16622 9288 19062 9344
rect 19118 9288 21086 9344
rect 21142 9288 21147 9344
rect 16622 9286 21147 9288
rect 19057 9283 19123 9286
rect 21081 9283 21147 9286
rect 25405 9346 25471 9349
rect 25957 9346 26023 9349
rect 25405 9344 26023 9346
rect 25405 9288 25410 9344
rect 25466 9288 25962 9344
rect 26018 9288 26023 9344
rect 25405 9286 26023 9288
rect 25405 9283 25471 9286
rect 25957 9283 26023 9286
rect 28758 9284 28764 9348
rect 28828 9346 28834 9348
rect 31385 9346 31451 9349
rect 28828 9344 31451 9346
rect 28828 9288 31390 9344
rect 31446 9288 31451 9344
rect 28828 9286 31451 9288
rect 28828 9284 28834 9286
rect 31385 9283 31451 9286
rect 5707 9280 6023 9281
rect 5707 9216 5713 9280
rect 5777 9216 5793 9280
rect 5857 9216 5873 9280
rect 5937 9216 5953 9280
rect 6017 9216 6023 9280
rect 5707 9215 6023 9216
rect 15229 9280 15545 9281
rect 15229 9216 15235 9280
rect 15299 9216 15315 9280
rect 15379 9216 15395 9280
rect 15459 9216 15475 9280
rect 15539 9216 15545 9280
rect 15229 9215 15545 9216
rect 24751 9280 25067 9281
rect 24751 9216 24757 9280
rect 24821 9216 24837 9280
rect 24901 9216 24917 9280
rect 24981 9216 24997 9280
rect 25061 9216 25067 9280
rect 24751 9215 25067 9216
rect 34273 9280 34589 9281
rect 34273 9216 34279 9280
rect 34343 9216 34359 9280
rect 34423 9216 34439 9280
rect 34503 9216 34519 9280
rect 34583 9216 34589 9280
rect 34273 9215 34589 9216
rect 10777 9210 10843 9213
rect 12525 9210 12591 9213
rect 10777 9208 12591 9210
rect 10777 9152 10782 9208
rect 10838 9152 12530 9208
rect 12586 9152 12591 9208
rect 10777 9150 12591 9152
rect 10777 9147 10843 9150
rect 12525 9147 12591 9150
rect 13169 9210 13235 9213
rect 13445 9210 13511 9213
rect 13169 9208 13511 9210
rect 13169 9152 13174 9208
rect 13230 9152 13450 9208
rect 13506 9152 13511 9208
rect 13169 9150 13511 9152
rect 13169 9147 13235 9150
rect 13445 9147 13511 9150
rect 16021 9210 16087 9213
rect 19517 9210 19583 9213
rect 25313 9210 25379 9213
rect 27889 9210 27955 9213
rect 30281 9210 30347 9213
rect 30414 9210 30420 9212
rect 16021 9208 24640 9210
rect 16021 9152 16026 9208
rect 16082 9152 19522 9208
rect 19578 9152 24640 9208
rect 16021 9150 24640 9152
rect 16021 9147 16087 9150
rect 19517 9147 19583 9150
rect 11881 9074 11947 9077
rect 14733 9074 14799 9077
rect 15101 9076 15167 9077
rect 11881 9072 14799 9074
rect 11881 9016 11886 9072
rect 11942 9016 14738 9072
rect 14794 9016 14799 9072
rect 11881 9014 14799 9016
rect 11881 9011 11947 9014
rect 14733 9011 14799 9014
rect 15096 9012 15102 9076
rect 15166 9074 15172 9076
rect 15377 9074 15443 9077
rect 20989 9074 21055 9077
rect 15166 9014 15254 9074
rect 15377 9072 21055 9074
rect 15377 9016 15382 9072
rect 15438 9016 20994 9072
rect 21050 9016 21055 9072
rect 15377 9014 21055 9016
rect 24580 9074 24640 9150
rect 25313 9208 26250 9210
rect 25313 9152 25318 9208
rect 25374 9152 26250 9208
rect 25313 9150 26250 9152
rect 25313 9147 25379 9150
rect 25957 9074 26023 9077
rect 24580 9072 26023 9074
rect 24580 9016 25962 9072
rect 26018 9016 26023 9072
rect 24580 9014 26023 9016
rect 26190 9074 26250 9150
rect 27889 9208 30420 9210
rect 27889 9152 27894 9208
rect 27950 9152 30286 9208
rect 30342 9152 30420 9208
rect 27889 9150 30420 9152
rect 27889 9147 27955 9150
rect 30281 9147 30347 9150
rect 30414 9148 30420 9150
rect 30484 9148 30490 9212
rect 31845 9210 31911 9213
rect 33685 9210 33751 9213
rect 31845 9208 33751 9210
rect 31845 9152 31850 9208
rect 31906 9152 33690 9208
rect 33746 9152 33751 9208
rect 31845 9150 33751 9152
rect 31845 9147 31911 9150
rect 33685 9147 33751 9150
rect 31017 9074 31083 9077
rect 26190 9072 31083 9074
rect 26190 9016 31022 9072
rect 31078 9016 31083 9072
rect 26190 9014 31083 9016
rect 15166 9012 15172 9014
rect 15101 9011 15167 9012
rect 15377 9011 15443 9014
rect 20989 9011 21055 9014
rect 25957 9011 26023 9014
rect 31017 9011 31083 9014
rect 31385 9074 31451 9077
rect 33317 9074 33383 9077
rect 31385 9072 33383 9074
rect 31385 9016 31390 9072
rect 31446 9016 33322 9072
rect 33378 9016 33383 9072
rect 31385 9014 33383 9016
rect 31385 9011 31451 9014
rect 33317 9011 33383 9014
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 9765 8938 9831 8941
rect 15929 8938 15995 8941
rect 18638 8938 18644 8940
rect 9765 8936 15995 8938
rect 9765 8880 9770 8936
rect 9826 8880 15934 8936
rect 15990 8880 15995 8936
rect 9765 8878 15995 8880
rect 9765 8875 9831 8878
rect 15929 8875 15995 8878
rect 16070 8878 18644 8938
rect 13169 8802 13235 8805
rect 16070 8802 16130 8878
rect 18638 8876 18644 8878
rect 18708 8876 18714 8940
rect 19333 8938 19399 8941
rect 19333 8936 24410 8938
rect 19333 8880 19338 8936
rect 19394 8880 24410 8936
rect 19333 8878 24410 8880
rect 19333 8875 19399 8878
rect 13169 8800 16130 8802
rect 13169 8744 13174 8800
rect 13230 8744 16130 8800
rect 13169 8742 16130 8744
rect 17309 8802 17375 8805
rect 19701 8802 19767 8805
rect 17309 8800 19767 8802
rect 17309 8744 17314 8800
rect 17370 8744 19706 8800
rect 19762 8744 19767 8800
rect 17309 8742 19767 8744
rect 13169 8739 13235 8742
rect 17309 8739 17375 8742
rect 19701 8739 19767 8742
rect 20662 8740 20668 8804
rect 20732 8802 20738 8804
rect 21909 8802 21975 8805
rect 20732 8800 21975 8802
rect 20732 8744 21914 8800
rect 21970 8744 21975 8800
rect 20732 8742 21975 8744
rect 24350 8802 24410 8878
rect 24526 8876 24532 8940
rect 24596 8938 24602 8940
rect 33777 8938 33843 8941
rect 24596 8936 33843 8938
rect 24596 8880 33782 8936
rect 33838 8880 33843 8936
rect 24596 8878 33843 8880
rect 24596 8876 24602 8878
rect 33777 8875 33843 8878
rect 34646 8876 34652 8940
rect 34716 8938 34722 8940
rect 36905 8938 36971 8941
rect 34716 8936 36971 8938
rect 34716 8880 36910 8936
rect 36966 8880 36971 8936
rect 34716 8878 36971 8880
rect 34716 8876 34722 8878
rect 36905 8875 36971 8878
rect 24669 8802 24735 8805
rect 28758 8802 28764 8804
rect 24350 8800 28764 8802
rect 24350 8744 24674 8800
rect 24730 8744 28764 8800
rect 24350 8742 28764 8744
rect 20732 8740 20738 8742
rect 21909 8739 21975 8742
rect 24669 8739 24735 8742
rect 28758 8740 28764 8742
rect 28828 8740 28834 8804
rect 31017 8802 31083 8805
rect 32121 8802 32187 8805
rect 32806 8802 32812 8804
rect 31017 8800 32812 8802
rect 31017 8744 31022 8800
rect 31078 8744 32126 8800
rect 32182 8744 32812 8800
rect 31017 8742 32812 8744
rect 31017 8739 31083 8742
rect 32121 8739 32187 8742
rect 32806 8740 32812 8742
rect 32876 8740 32882 8804
rect 32990 8740 32996 8804
rect 33060 8802 33066 8804
rect 34605 8802 34671 8805
rect 33060 8800 34671 8802
rect 33060 8744 34610 8800
rect 34666 8744 34671 8800
rect 33060 8742 34671 8744
rect 33060 8740 33066 8742
rect 34605 8739 34671 8742
rect 10468 8736 10784 8737
rect 10468 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10784 8736
rect 10468 8671 10784 8672
rect 19990 8736 20306 8737
rect 19990 8672 19996 8736
rect 20060 8672 20076 8736
rect 20140 8672 20156 8736
rect 20220 8672 20236 8736
rect 20300 8672 20306 8736
rect 19990 8671 20306 8672
rect 29512 8736 29828 8737
rect 29512 8672 29518 8736
rect 29582 8672 29598 8736
rect 29662 8672 29678 8736
rect 29742 8672 29758 8736
rect 29822 8672 29828 8736
rect 29512 8671 29828 8672
rect 39034 8736 39350 8737
rect 39034 8672 39040 8736
rect 39104 8672 39120 8736
rect 39184 8672 39200 8736
rect 39264 8672 39280 8736
rect 39344 8672 39350 8736
rect 39034 8671 39350 8672
rect 4061 8666 4127 8669
rect 4613 8666 4679 8669
rect 4061 8664 4679 8666
rect 4061 8608 4066 8664
rect 4122 8608 4618 8664
rect 4674 8608 4679 8664
rect 4061 8606 4679 8608
rect 4061 8603 4127 8606
rect 4613 8603 4679 8606
rect 7005 8668 7071 8669
rect 7005 8664 7052 8668
rect 7116 8666 7122 8668
rect 11145 8666 11211 8669
rect 17493 8666 17559 8669
rect 20989 8666 21055 8669
rect 28073 8666 28139 8669
rect 28390 8666 28396 8668
rect 7005 8608 7010 8664
rect 7005 8604 7052 8608
rect 7116 8606 7162 8666
rect 11145 8664 17602 8666
rect 11145 8608 11150 8664
rect 11206 8608 17498 8664
rect 17554 8608 17602 8664
rect 11145 8606 17602 8608
rect 7116 8604 7122 8606
rect 7005 8603 7071 8604
rect 11145 8603 11211 8606
rect 17493 8603 17602 8606
rect 20989 8664 26986 8666
rect 20989 8608 20994 8664
rect 21050 8608 26986 8664
rect 20989 8606 26986 8608
rect 20989 8603 21055 8606
rect 3417 8530 3483 8533
rect 5441 8530 5507 8533
rect 7097 8530 7163 8533
rect 7649 8530 7715 8533
rect 17542 8530 17602 8603
rect 20989 8530 21055 8533
rect 3417 8528 7715 8530
rect 3417 8472 3422 8528
rect 3478 8472 5446 8528
rect 5502 8472 7102 8528
rect 7158 8472 7654 8528
rect 7710 8472 7715 8528
rect 3417 8470 7715 8472
rect 3417 8467 3483 8470
rect 5441 8467 5507 8470
rect 7097 8467 7163 8470
rect 7649 8467 7715 8470
rect 10182 8470 17234 8530
rect 17542 8528 21055 8530
rect 17542 8472 20994 8528
rect 21050 8472 21055 8528
rect 17542 8470 21055 8472
rect 10182 8397 10242 8470
rect 6453 8394 6519 8397
rect 10133 8394 10242 8397
rect 6453 8392 10242 8394
rect 6453 8336 6458 8392
rect 6514 8336 10138 8392
rect 10194 8336 10242 8392
rect 6453 8334 10242 8336
rect 10777 8394 10843 8397
rect 17033 8394 17099 8397
rect 10777 8392 17099 8394
rect 10777 8336 10782 8392
rect 10838 8336 17038 8392
rect 17094 8336 17099 8392
rect 10777 8334 17099 8336
rect 17174 8394 17234 8470
rect 20989 8467 21055 8470
rect 21449 8530 21515 8533
rect 25589 8530 25655 8533
rect 26182 8530 26188 8532
rect 21449 8528 25330 8530
rect 21449 8472 21454 8528
rect 21510 8472 25330 8528
rect 21449 8470 25330 8472
rect 21449 8467 21515 8470
rect 22185 8394 22251 8397
rect 17174 8392 22251 8394
rect 17174 8336 22190 8392
rect 22246 8336 22251 8392
rect 17174 8334 22251 8336
rect 6453 8331 6519 8334
rect 10133 8331 10199 8334
rect 10777 8331 10843 8334
rect 17033 8331 17099 8334
rect 22185 8331 22251 8334
rect 22369 8394 22435 8397
rect 25270 8394 25330 8470
rect 25589 8528 26188 8530
rect 25589 8472 25594 8528
rect 25650 8472 26188 8528
rect 25589 8470 26188 8472
rect 25589 8467 25655 8470
rect 26182 8468 26188 8470
rect 26252 8468 26258 8532
rect 26926 8530 26986 8606
rect 28073 8664 28396 8666
rect 28073 8608 28078 8664
rect 28134 8608 28396 8664
rect 28073 8606 28396 8608
rect 28073 8603 28139 8606
rect 28390 8604 28396 8606
rect 28460 8604 28466 8668
rect 28574 8604 28580 8668
rect 28644 8666 28650 8668
rect 28901 8666 28967 8669
rect 28644 8664 28967 8666
rect 28644 8608 28906 8664
rect 28962 8608 28967 8664
rect 28644 8606 28967 8608
rect 28644 8604 28650 8606
rect 28901 8603 28967 8606
rect 30281 8666 30347 8669
rect 34973 8666 35039 8669
rect 30281 8664 35039 8666
rect 30281 8608 30286 8664
rect 30342 8608 34978 8664
rect 35034 8608 35039 8664
rect 30281 8606 35039 8608
rect 30281 8603 30347 8606
rect 34973 8603 35039 8606
rect 37365 8530 37431 8533
rect 26926 8528 37431 8530
rect 26926 8472 37370 8528
rect 37426 8472 37431 8528
rect 26926 8470 37431 8472
rect 37365 8467 37431 8470
rect 27981 8394 28047 8397
rect 30557 8394 30623 8397
rect 22369 8392 25192 8394
rect 22369 8336 22374 8392
rect 22430 8336 25192 8392
rect 22369 8334 25192 8336
rect 25270 8392 30623 8394
rect 25270 8336 27986 8392
rect 28042 8336 30562 8392
rect 30618 8336 30623 8392
rect 25270 8334 30623 8336
rect 22369 8331 22435 8334
rect 6870 8198 9322 8258
rect 5707 8192 6023 8193
rect 5707 8128 5713 8192
rect 5777 8128 5793 8192
rect 5857 8128 5873 8192
rect 5937 8128 5953 8192
rect 6017 8128 6023 8192
rect 5707 8127 6023 8128
rect 2773 7986 2839 7989
rect 2773 7984 2882 7986
rect 2773 7928 2778 7984
rect 2834 7928 2882 7984
rect 2773 7923 2882 7928
rect 3182 7924 3188 7988
rect 3252 7986 3258 7988
rect 6870 7986 6930 8198
rect 9262 8122 9322 8198
rect 9438 8196 9444 8260
rect 9508 8258 9514 8260
rect 11605 8258 11671 8261
rect 21357 8258 21423 8261
rect 9508 8256 11671 8258
rect 9508 8200 11610 8256
rect 11666 8200 11671 8256
rect 9508 8198 11671 8200
rect 9508 8196 9514 8198
rect 11605 8195 11671 8198
rect 15656 8256 21423 8258
rect 15656 8200 21362 8256
rect 21418 8200 21423 8256
rect 15656 8198 21423 8200
rect 15229 8192 15545 8193
rect 15229 8128 15235 8192
rect 15299 8128 15315 8192
rect 15379 8128 15395 8192
rect 15459 8128 15475 8192
rect 15539 8128 15545 8192
rect 15229 8127 15545 8128
rect 11237 8122 11303 8125
rect 13486 8122 13492 8124
rect 9262 8120 11303 8122
rect 9262 8064 11242 8120
rect 11298 8064 11303 8120
rect 9262 8062 11303 8064
rect 11237 8059 11303 8062
rect 11470 8062 13492 8122
rect 3252 7926 6930 7986
rect 7649 7986 7715 7989
rect 10317 7986 10383 7989
rect 7649 7984 10383 7986
rect 7649 7928 7654 7984
rect 7710 7928 10322 7984
rect 10378 7928 10383 7984
rect 7649 7926 10383 7928
rect 3252 7924 3258 7926
rect 7649 7923 7715 7926
rect 10317 7923 10383 7926
rect 10685 7986 10751 7989
rect 11470 7986 11530 8062
rect 13486 8060 13492 8062
rect 13556 8060 13562 8124
rect 14365 8122 14431 8125
rect 15101 8122 15167 8125
rect 14365 8120 15167 8122
rect 14365 8064 14370 8120
rect 14426 8064 15106 8120
rect 15162 8064 15167 8120
rect 14365 8062 15167 8064
rect 14365 8059 14431 8062
rect 15101 8059 15167 8062
rect 10685 7984 11530 7986
rect 10685 7928 10690 7984
rect 10746 7928 11530 7984
rect 10685 7926 11530 7928
rect 12065 7986 12131 7989
rect 15656 7986 15716 8198
rect 21357 8195 21423 8198
rect 24751 8192 25067 8193
rect 24751 8128 24757 8192
rect 24821 8128 24837 8192
rect 24901 8128 24917 8192
rect 24981 8128 24997 8192
rect 25061 8128 25067 8192
rect 24751 8127 25067 8128
rect 17217 8122 17283 8125
rect 23289 8122 23355 8125
rect 17217 8120 23355 8122
rect 17217 8064 17222 8120
rect 17278 8064 23294 8120
rect 23350 8064 23355 8120
rect 17217 8062 23355 8064
rect 25132 8122 25192 8334
rect 27981 8331 28047 8334
rect 30557 8331 30623 8334
rect 31201 8394 31267 8397
rect 33041 8394 33107 8397
rect 38193 8394 38259 8397
rect 31201 8392 33107 8394
rect 31201 8336 31206 8392
rect 31262 8336 33046 8392
rect 33102 8336 33107 8392
rect 31201 8334 33107 8336
rect 31201 8331 31267 8334
rect 33041 8331 33107 8334
rect 33320 8392 38259 8394
rect 33320 8336 38198 8392
rect 38254 8336 38259 8392
rect 33320 8334 38259 8336
rect 31293 8258 31359 8261
rect 27662 8256 31359 8258
rect 27662 8200 31298 8256
rect 31354 8200 31359 8256
rect 27662 8198 31359 8200
rect 27662 8122 27722 8198
rect 31293 8195 31359 8198
rect 32949 8258 33015 8261
rect 33320 8258 33380 8334
rect 38193 8331 38259 8334
rect 32949 8256 33380 8258
rect 32949 8200 32954 8256
rect 33010 8200 33380 8256
rect 32949 8198 33380 8200
rect 32949 8195 33015 8198
rect 34273 8192 34589 8193
rect 34273 8128 34279 8192
rect 34343 8128 34359 8192
rect 34423 8128 34439 8192
rect 34503 8128 34519 8192
rect 34583 8128 34589 8192
rect 34273 8127 34589 8128
rect 25132 8062 27722 8122
rect 28625 8122 28691 8125
rect 28809 8122 28875 8125
rect 28625 8120 28875 8122
rect 28625 8064 28630 8120
rect 28686 8064 28814 8120
rect 28870 8064 28875 8120
rect 28625 8062 28875 8064
rect 17217 8059 17283 8062
rect 23289 8059 23355 8062
rect 28625 8059 28691 8062
rect 28809 8059 28875 8062
rect 29126 8060 29132 8124
rect 29196 8122 29202 8124
rect 29361 8122 29427 8125
rect 29196 8120 29427 8122
rect 29196 8064 29366 8120
rect 29422 8064 29427 8120
rect 29196 8062 29427 8064
rect 29196 8060 29202 8062
rect 29361 8059 29427 8062
rect 29821 8122 29887 8125
rect 33501 8122 33567 8125
rect 33685 8122 33751 8125
rect 29821 8120 33426 8122
rect 29821 8064 29826 8120
rect 29882 8064 33426 8120
rect 29821 8062 33426 8064
rect 29821 8059 29887 8062
rect 12065 7984 15716 7986
rect 12065 7928 12070 7984
rect 12126 7928 15716 7984
rect 12065 7926 15716 7928
rect 16757 7986 16823 7989
rect 24526 7986 24532 7988
rect 16757 7984 24532 7986
rect 16757 7928 16762 7984
rect 16818 7928 24532 7984
rect 16757 7926 24532 7928
rect 10685 7923 10751 7926
rect 12065 7923 12131 7926
rect 16757 7923 16823 7926
rect 24526 7924 24532 7926
rect 24596 7924 24602 7988
rect 24761 7986 24827 7989
rect 26049 7986 26115 7989
rect 24761 7984 26115 7986
rect 24761 7928 24766 7984
rect 24822 7928 26054 7984
rect 26110 7928 26115 7984
rect 24761 7926 26115 7928
rect 24761 7923 24827 7926
rect 26049 7923 26115 7926
rect 28073 7986 28139 7989
rect 30281 7986 30347 7989
rect 28073 7984 30347 7986
rect 28073 7928 28078 7984
rect 28134 7928 30286 7984
rect 30342 7928 30347 7984
rect 28073 7926 30347 7928
rect 33366 7986 33426 8062
rect 33501 8120 33751 8122
rect 33501 8064 33506 8120
rect 33562 8064 33690 8120
rect 33746 8064 33751 8120
rect 33501 8062 33751 8064
rect 33501 8059 33567 8062
rect 33685 8059 33751 8062
rect 34697 8122 34763 8125
rect 37549 8122 37615 8125
rect 37733 8122 37799 8125
rect 34697 8120 37799 8122
rect 34697 8064 34702 8120
rect 34758 8064 37554 8120
rect 37610 8064 37738 8120
rect 37794 8064 37799 8120
rect 34697 8062 37799 8064
rect 34697 8059 34763 8062
rect 37549 8059 37615 8062
rect 37733 8059 37799 8062
rect 37733 7986 37799 7989
rect 33366 7984 37799 7986
rect 33366 7928 37738 7984
rect 37794 7928 37799 7984
rect 33366 7926 37799 7928
rect 28073 7923 28139 7926
rect 30281 7923 30347 7926
rect 37733 7923 37799 7926
rect 0 7578 800 7608
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 2822 7173 2882 7923
rect 9857 7850 9923 7853
rect 18781 7850 18847 7853
rect 9857 7848 18847 7850
rect 9857 7792 9862 7848
rect 9918 7792 18786 7848
rect 18842 7792 18847 7848
rect 9857 7790 18847 7792
rect 9857 7787 9923 7790
rect 18781 7787 18847 7790
rect 19701 7850 19767 7853
rect 36261 7850 36327 7853
rect 19701 7848 36327 7850
rect 19701 7792 19706 7848
rect 19762 7792 36266 7848
rect 36322 7792 36327 7848
rect 19701 7790 36327 7792
rect 19701 7787 19767 7790
rect 36261 7787 36327 7790
rect 3601 7714 3667 7717
rect 8017 7714 8083 7717
rect 3601 7712 8083 7714
rect 3601 7656 3606 7712
rect 3662 7656 8022 7712
rect 8078 7656 8083 7712
rect 3601 7654 8083 7656
rect 3601 7651 3667 7654
rect 8017 7651 8083 7654
rect 12249 7714 12315 7717
rect 17493 7714 17559 7717
rect 12249 7712 17559 7714
rect 12249 7656 12254 7712
rect 12310 7656 17498 7712
rect 17554 7656 17559 7712
rect 12249 7654 17559 7656
rect 12249 7651 12315 7654
rect 17493 7651 17559 7654
rect 20529 7714 20595 7717
rect 22277 7714 22343 7717
rect 20529 7712 22343 7714
rect 20529 7656 20534 7712
rect 20590 7656 22282 7712
rect 22338 7656 22343 7712
rect 20529 7654 22343 7656
rect 20529 7651 20595 7654
rect 22277 7651 22343 7654
rect 23422 7652 23428 7716
rect 23492 7714 23498 7716
rect 26049 7714 26115 7717
rect 23492 7712 26115 7714
rect 23492 7656 26054 7712
rect 26110 7656 26115 7712
rect 23492 7654 26115 7656
rect 23492 7652 23498 7654
rect 26049 7651 26115 7654
rect 26417 7714 26483 7717
rect 28901 7714 28967 7717
rect 26417 7712 28967 7714
rect 26417 7656 26422 7712
rect 26478 7656 28906 7712
rect 28962 7656 28967 7712
rect 26417 7654 28967 7656
rect 26417 7651 26483 7654
rect 28901 7651 28967 7654
rect 30557 7714 30623 7717
rect 30925 7714 30991 7717
rect 37181 7714 37247 7717
rect 30557 7712 37247 7714
rect 30557 7656 30562 7712
rect 30618 7656 30930 7712
rect 30986 7656 37186 7712
rect 37242 7656 37247 7712
rect 30557 7654 37247 7656
rect 30557 7651 30623 7654
rect 30925 7651 30991 7654
rect 37181 7651 37247 7654
rect 10468 7648 10784 7649
rect 10468 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10784 7648
rect 10468 7583 10784 7584
rect 19990 7648 20306 7649
rect 19990 7584 19996 7648
rect 20060 7584 20076 7648
rect 20140 7584 20156 7648
rect 20220 7584 20236 7648
rect 20300 7584 20306 7648
rect 19990 7583 20306 7584
rect 29512 7648 29828 7649
rect 29512 7584 29518 7648
rect 29582 7584 29598 7648
rect 29662 7584 29678 7648
rect 29742 7584 29758 7648
rect 29822 7584 29828 7648
rect 29512 7583 29828 7584
rect 39034 7648 39350 7649
rect 39034 7584 39040 7648
rect 39104 7584 39120 7648
rect 39184 7584 39200 7648
rect 39264 7584 39280 7648
rect 39344 7584 39350 7648
rect 39034 7583 39350 7584
rect 4061 7578 4127 7581
rect 5717 7578 5783 7581
rect 8109 7578 8175 7581
rect 4061 7576 8175 7578
rect 4061 7520 4066 7576
rect 4122 7520 5722 7576
rect 5778 7520 8114 7576
rect 8170 7520 8175 7576
rect 4061 7518 8175 7520
rect 4061 7515 4127 7518
rect 5717 7515 5783 7518
rect 8109 7515 8175 7518
rect 11237 7578 11303 7581
rect 16941 7578 17007 7581
rect 17309 7578 17375 7581
rect 27061 7578 27127 7581
rect 27705 7578 27771 7581
rect 11237 7576 19810 7578
rect 11237 7520 11242 7576
rect 11298 7520 16946 7576
rect 17002 7520 17314 7576
rect 17370 7520 19810 7576
rect 11237 7518 19810 7520
rect 11237 7515 11303 7518
rect 16941 7515 17007 7518
rect 17309 7515 17375 7518
rect 4797 7442 4863 7445
rect 17217 7442 17283 7445
rect 4797 7440 17283 7442
rect 4797 7384 4802 7440
rect 4858 7384 17222 7440
rect 17278 7384 17283 7440
rect 4797 7382 17283 7384
rect 19750 7442 19810 7518
rect 24902 7576 27771 7578
rect 24902 7520 27066 7576
rect 27122 7520 27710 7576
rect 27766 7520 27771 7576
rect 24902 7518 27771 7520
rect 23749 7442 23815 7445
rect 19750 7440 23815 7442
rect 19750 7384 23754 7440
rect 23810 7384 23815 7440
rect 19750 7382 23815 7384
rect 4797 7379 4863 7382
rect 17217 7379 17283 7382
rect 23749 7379 23815 7382
rect 4337 7306 4403 7309
rect 4889 7306 4955 7309
rect 5809 7306 5875 7309
rect 4337 7304 5875 7306
rect 4337 7248 4342 7304
rect 4398 7248 4894 7304
rect 4950 7248 5814 7304
rect 5870 7248 5875 7304
rect 4337 7246 5875 7248
rect 4337 7243 4403 7246
rect 4889 7243 4955 7246
rect 5809 7243 5875 7246
rect 8937 7306 9003 7309
rect 21449 7306 21515 7309
rect 23841 7306 23907 7309
rect 24902 7306 24962 7518
rect 27061 7515 27127 7518
rect 27705 7515 27771 7518
rect 29913 7578 29979 7581
rect 35157 7578 35223 7581
rect 39566 7578 40366 7608
rect 29913 7576 35223 7578
rect 29913 7520 29918 7576
rect 29974 7520 35162 7576
rect 35218 7520 35223 7576
rect 29913 7518 35223 7520
rect 29913 7515 29979 7518
rect 35157 7515 35223 7518
rect 39438 7518 40366 7578
rect 25037 7442 25103 7445
rect 25313 7442 25379 7445
rect 25037 7440 25379 7442
rect 25037 7384 25042 7440
rect 25098 7384 25318 7440
rect 25374 7384 25379 7440
rect 25037 7382 25379 7384
rect 25037 7379 25103 7382
rect 25313 7379 25379 7382
rect 25497 7442 25563 7445
rect 32673 7442 32739 7445
rect 25497 7440 32739 7442
rect 25497 7384 25502 7440
rect 25558 7384 32678 7440
rect 32734 7384 32739 7440
rect 25497 7382 32739 7384
rect 25497 7379 25563 7382
rect 32673 7379 32739 7382
rect 38653 7442 38719 7445
rect 39438 7442 39498 7518
rect 39566 7488 40366 7518
rect 38653 7440 39498 7442
rect 38653 7384 38658 7440
rect 38714 7384 39498 7440
rect 38653 7382 39498 7384
rect 38653 7379 38719 7382
rect 8937 7304 21515 7306
rect 8937 7248 8942 7304
rect 8998 7248 21454 7304
rect 21510 7248 21515 7304
rect 8937 7246 21515 7248
rect 8937 7243 9003 7246
rect 21449 7243 21515 7246
rect 21590 7304 24962 7306
rect 21590 7248 23846 7304
rect 23902 7248 24962 7304
rect 21590 7246 24962 7248
rect 25221 7306 25287 7309
rect 29913 7306 29979 7309
rect 36077 7306 36143 7309
rect 25221 7304 29979 7306
rect 25221 7248 25226 7304
rect 25282 7248 29918 7304
rect 29974 7248 29979 7304
rect 25221 7246 29979 7248
rect 2773 7168 2882 7173
rect 2773 7112 2778 7168
rect 2834 7112 2882 7168
rect 2773 7110 2882 7112
rect 10317 7170 10383 7173
rect 10501 7170 10567 7173
rect 14917 7170 14983 7173
rect 10317 7168 14983 7170
rect 10317 7112 10322 7168
rect 10378 7112 10506 7168
rect 10562 7112 14922 7168
rect 14978 7112 14983 7168
rect 10317 7110 14983 7112
rect 2773 7107 2839 7110
rect 10317 7107 10383 7110
rect 10501 7107 10567 7110
rect 14917 7107 14983 7110
rect 15745 7170 15811 7173
rect 21590 7170 21650 7246
rect 23841 7243 23907 7246
rect 25221 7243 25287 7246
rect 29913 7243 29979 7246
rect 31710 7304 36143 7306
rect 31710 7248 36082 7304
rect 36138 7248 36143 7304
rect 31710 7246 36143 7248
rect 15745 7168 21650 7170
rect 15745 7112 15750 7168
rect 15806 7112 21650 7168
rect 15745 7110 21650 7112
rect 25313 7170 25379 7173
rect 31710 7170 31770 7246
rect 36077 7243 36143 7246
rect 25313 7168 31770 7170
rect 25313 7112 25318 7168
rect 25374 7112 31770 7168
rect 25313 7110 31770 7112
rect 15745 7107 15811 7110
rect 25313 7107 25379 7110
rect 5707 7104 6023 7105
rect 5707 7040 5713 7104
rect 5777 7040 5793 7104
rect 5857 7040 5873 7104
rect 5937 7040 5953 7104
rect 6017 7040 6023 7104
rect 5707 7039 6023 7040
rect 15229 7104 15545 7105
rect 15229 7040 15235 7104
rect 15299 7040 15315 7104
rect 15379 7040 15395 7104
rect 15459 7040 15475 7104
rect 15539 7040 15545 7104
rect 15229 7039 15545 7040
rect 24751 7104 25067 7105
rect 24751 7040 24757 7104
rect 24821 7040 24837 7104
rect 24901 7040 24917 7104
rect 24981 7040 24997 7104
rect 25061 7040 25067 7104
rect 24751 7039 25067 7040
rect 34273 7104 34589 7105
rect 34273 7040 34279 7104
rect 34343 7040 34359 7104
rect 34423 7040 34439 7104
rect 34503 7040 34519 7104
rect 34583 7040 34589 7104
rect 34273 7039 34589 7040
rect 12433 7034 12499 7037
rect 12566 7034 12572 7036
rect 12433 7032 12572 7034
rect 12433 6976 12438 7032
rect 12494 6976 12572 7032
rect 12433 6974 12572 6976
rect 12433 6971 12499 6974
rect 12566 6972 12572 6974
rect 12636 6972 12642 7036
rect 16389 7034 16455 7037
rect 17585 7034 17651 7037
rect 16389 7032 17651 7034
rect 16389 6976 16394 7032
rect 16450 6976 17590 7032
rect 17646 6976 17651 7032
rect 16389 6974 17651 6976
rect 16389 6971 16455 6974
rect 17585 6971 17651 6974
rect 19793 7034 19859 7037
rect 22001 7034 22067 7037
rect 19793 7032 22067 7034
rect 19793 6976 19798 7032
rect 19854 6976 22006 7032
rect 22062 6976 22067 7032
rect 19793 6974 22067 6976
rect 19793 6971 19859 6974
rect 22001 6971 22067 6974
rect 22737 7034 22803 7037
rect 25221 7034 25287 7037
rect 31017 7034 31083 7037
rect 22737 7032 24594 7034
rect 22737 6976 22742 7032
rect 22798 6976 24594 7032
rect 22737 6974 24594 6976
rect 22737 6971 22803 6974
rect 3049 6898 3115 6901
rect 4102 6898 4108 6900
rect 3049 6896 4108 6898
rect 3049 6840 3054 6896
rect 3110 6840 4108 6896
rect 3049 6838 4108 6840
rect 3049 6835 3115 6838
rect 4102 6836 4108 6838
rect 4172 6836 4178 6900
rect 4521 6898 4587 6901
rect 7281 6898 7347 6901
rect 4521 6896 7347 6898
rect 4521 6840 4526 6896
rect 4582 6840 7286 6896
rect 7342 6840 7347 6896
rect 4521 6838 7347 6840
rect 4521 6835 4587 6838
rect 7281 6835 7347 6838
rect 10869 6898 10935 6901
rect 20805 6898 20871 6901
rect 24301 6898 24367 6901
rect 10869 6896 24367 6898
rect 10869 6840 10874 6896
rect 10930 6840 20810 6896
rect 20866 6840 24306 6896
rect 24362 6840 24367 6896
rect 10869 6838 24367 6840
rect 24534 6898 24594 6974
rect 25221 7032 31083 7034
rect 25221 6976 25226 7032
rect 25282 6976 31022 7032
rect 31078 6976 31083 7032
rect 25221 6974 31083 6976
rect 25221 6971 25287 6974
rect 31017 6971 31083 6974
rect 31201 7034 31267 7037
rect 32857 7034 32923 7037
rect 31201 7032 32923 7034
rect 31201 6976 31206 7032
rect 31262 6976 32862 7032
rect 32918 6976 32923 7032
rect 31201 6974 32923 6976
rect 31201 6971 31267 6974
rect 32857 6971 32923 6974
rect 26693 6898 26759 6901
rect 24534 6896 26759 6898
rect 24534 6840 26698 6896
rect 26754 6840 26759 6896
rect 24534 6838 26759 6840
rect 10869 6835 10935 6838
rect 20805 6835 20871 6838
rect 24301 6835 24367 6838
rect 26693 6835 26759 6838
rect 27705 6898 27771 6901
rect 30005 6898 30071 6901
rect 27705 6896 30071 6898
rect 27705 6840 27710 6896
rect 27766 6840 30010 6896
rect 30066 6840 30071 6896
rect 27705 6838 30071 6840
rect 27705 6835 27771 6838
rect 30005 6835 30071 6838
rect 30925 6898 30991 6901
rect 31150 6898 31156 6900
rect 30925 6896 31156 6898
rect 30925 6840 30930 6896
rect 30986 6840 31156 6896
rect 30925 6838 31156 6840
rect 30925 6835 30991 6838
rect 31150 6836 31156 6838
rect 31220 6836 31226 6900
rect 33501 6898 33567 6901
rect 34237 6898 34303 6901
rect 33501 6896 34303 6898
rect 33501 6840 33506 6896
rect 33562 6840 34242 6896
rect 34298 6840 34303 6896
rect 33501 6838 34303 6840
rect 33501 6835 33567 6838
rect 34237 6835 34303 6838
rect 6453 6764 6519 6765
rect 6453 6760 6500 6764
rect 6564 6762 6570 6764
rect 6913 6762 6979 6765
rect 7046 6762 7052 6764
rect 6453 6704 6458 6760
rect 6453 6700 6500 6704
rect 6564 6702 6610 6762
rect 6913 6760 7052 6762
rect 6913 6704 6918 6760
rect 6974 6704 7052 6760
rect 6913 6702 7052 6704
rect 6564 6700 6570 6702
rect 6453 6699 6519 6700
rect 6913 6699 6979 6702
rect 7046 6700 7052 6702
rect 7116 6700 7122 6764
rect 9622 6700 9628 6764
rect 9692 6762 9698 6764
rect 12525 6762 12591 6765
rect 15694 6762 15700 6764
rect 9692 6702 12450 6762
rect 9692 6700 9698 6702
rect 5349 6626 5415 6629
rect 7189 6626 7255 6629
rect 5349 6624 7255 6626
rect 5349 6568 5354 6624
rect 5410 6568 7194 6624
rect 7250 6568 7255 6624
rect 5349 6566 7255 6568
rect 12390 6626 12450 6702
rect 12525 6760 15700 6762
rect 12525 6704 12530 6760
rect 12586 6704 15700 6760
rect 12525 6702 15700 6704
rect 12525 6699 12591 6702
rect 15694 6700 15700 6702
rect 15764 6700 15770 6764
rect 15837 6762 15903 6765
rect 25313 6762 25379 6765
rect 34881 6762 34947 6765
rect 15837 6760 25379 6762
rect 15837 6704 15842 6760
rect 15898 6704 25318 6760
rect 25374 6704 25379 6760
rect 15837 6702 25379 6704
rect 15837 6699 15903 6702
rect 25313 6699 25379 6702
rect 28030 6760 34947 6762
rect 28030 6704 34886 6760
rect 34942 6704 34947 6760
rect 28030 6702 34947 6704
rect 17953 6626 18019 6629
rect 22369 6628 22435 6629
rect 22318 6626 22324 6628
rect 12390 6624 18019 6626
rect 12390 6568 17958 6624
rect 18014 6568 18019 6624
rect 12390 6566 18019 6568
rect 22278 6566 22324 6626
rect 22388 6624 22435 6628
rect 22430 6568 22435 6624
rect 5349 6563 5415 6566
rect 7189 6563 7255 6566
rect 17953 6563 18019 6566
rect 22318 6564 22324 6566
rect 22388 6564 22435 6568
rect 22369 6563 22435 6564
rect 24117 6626 24183 6629
rect 28030 6626 28090 6702
rect 34881 6699 34947 6702
rect 35249 6762 35315 6765
rect 36905 6762 36971 6765
rect 35249 6760 36971 6762
rect 35249 6704 35254 6760
rect 35310 6704 36910 6760
rect 36966 6704 36971 6760
rect 35249 6702 36971 6704
rect 35249 6699 35315 6702
rect 36905 6699 36971 6702
rect 24117 6624 28090 6626
rect 24117 6568 24122 6624
rect 24178 6568 28090 6624
rect 24117 6566 28090 6568
rect 34053 6626 34119 6629
rect 36077 6626 36143 6629
rect 34053 6624 36143 6626
rect 34053 6568 34058 6624
rect 34114 6568 36082 6624
rect 36138 6568 36143 6624
rect 34053 6566 36143 6568
rect 24117 6563 24183 6566
rect 34053 6563 34119 6566
rect 36077 6563 36143 6566
rect 10468 6560 10784 6561
rect 10468 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10784 6560
rect 10468 6495 10784 6496
rect 19990 6560 20306 6561
rect 19990 6496 19996 6560
rect 20060 6496 20076 6560
rect 20140 6496 20156 6560
rect 20220 6496 20236 6560
rect 20300 6496 20306 6560
rect 19990 6495 20306 6496
rect 29512 6560 29828 6561
rect 29512 6496 29518 6560
rect 29582 6496 29598 6560
rect 29662 6496 29678 6560
rect 29742 6496 29758 6560
rect 29822 6496 29828 6560
rect 29512 6495 29828 6496
rect 39034 6560 39350 6561
rect 39034 6496 39040 6560
rect 39104 6496 39120 6560
rect 39184 6496 39200 6560
rect 39264 6496 39280 6560
rect 39344 6496 39350 6560
rect 39034 6495 39350 6496
rect 3141 6490 3207 6493
rect 3509 6490 3575 6493
rect 9213 6490 9279 6493
rect 9857 6490 9923 6493
rect 3141 6488 8218 6490
rect 3141 6432 3146 6488
rect 3202 6432 3514 6488
rect 3570 6432 8218 6488
rect 3141 6430 8218 6432
rect 3141 6427 3207 6430
rect 3509 6427 3575 6430
rect 5165 6354 5231 6357
rect 8017 6354 8083 6357
rect 5165 6352 8083 6354
rect 5165 6296 5170 6352
rect 5226 6296 8022 6352
rect 8078 6296 8083 6352
rect 5165 6294 8083 6296
rect 8158 6354 8218 6430
rect 9213 6488 9923 6490
rect 9213 6432 9218 6488
rect 9274 6432 9862 6488
rect 9918 6432 9923 6488
rect 9213 6430 9923 6432
rect 9213 6427 9279 6430
rect 9857 6427 9923 6430
rect 13537 6490 13603 6493
rect 13854 6490 13860 6492
rect 13537 6488 13860 6490
rect 13537 6432 13542 6488
rect 13598 6432 13860 6488
rect 13537 6430 13860 6432
rect 13537 6427 13603 6430
rect 13854 6428 13860 6430
rect 13924 6428 13930 6492
rect 14549 6490 14615 6493
rect 16481 6490 16547 6493
rect 17493 6490 17559 6493
rect 14549 6488 17559 6490
rect 14549 6432 14554 6488
rect 14610 6432 16486 6488
rect 16542 6432 17498 6488
rect 17554 6432 17559 6488
rect 14549 6430 17559 6432
rect 14549 6427 14615 6430
rect 16481 6427 16547 6430
rect 17493 6427 17559 6430
rect 20529 6490 20595 6493
rect 26918 6490 26924 6492
rect 20529 6488 26924 6490
rect 20529 6432 20534 6488
rect 20590 6432 26924 6488
rect 20529 6430 26924 6432
rect 20529 6427 20595 6430
rect 26918 6428 26924 6430
rect 26988 6490 26994 6492
rect 30005 6490 30071 6493
rect 32673 6490 32739 6493
rect 35893 6490 35959 6493
rect 26988 6430 29010 6490
rect 26988 6428 26994 6430
rect 10041 6354 10107 6357
rect 10501 6354 10567 6357
rect 8158 6294 9920 6354
rect 5165 6291 5231 6294
rect 8017 6291 8083 6294
rect 9581 6218 9647 6221
rect 3558 6216 9647 6218
rect 3558 6160 9586 6216
rect 9642 6160 9647 6216
rect 3558 6158 9647 6160
rect 9860 6218 9920 6294
rect 10041 6352 10567 6354
rect 10041 6296 10046 6352
rect 10102 6296 10506 6352
rect 10562 6296 10567 6352
rect 10041 6294 10567 6296
rect 10041 6291 10107 6294
rect 10501 6291 10567 6294
rect 11053 6354 11119 6357
rect 16573 6354 16639 6357
rect 11053 6352 16639 6354
rect 11053 6296 11058 6352
rect 11114 6296 16578 6352
rect 16634 6296 16639 6352
rect 11053 6294 16639 6296
rect 11053 6291 11119 6294
rect 16573 6291 16639 6294
rect 19558 6292 19564 6356
rect 19628 6354 19634 6356
rect 20437 6354 20503 6357
rect 19628 6352 20503 6354
rect 19628 6296 20442 6352
rect 20498 6296 20503 6352
rect 19628 6294 20503 6296
rect 19628 6292 19634 6294
rect 20437 6291 20503 6294
rect 20621 6354 20687 6357
rect 22461 6354 22527 6357
rect 25814 6354 25820 6356
rect 20621 6352 22110 6354
rect 20621 6296 20626 6352
rect 20682 6296 22110 6352
rect 20621 6294 22110 6296
rect 20621 6291 20687 6294
rect 12525 6218 12591 6221
rect 22050 6218 22110 6294
rect 22461 6352 25820 6354
rect 22461 6296 22466 6352
rect 22522 6296 25820 6352
rect 22461 6294 25820 6296
rect 22461 6291 22527 6294
rect 25814 6292 25820 6294
rect 25884 6292 25890 6356
rect 28950 6354 29010 6430
rect 30005 6488 30666 6490
rect 30005 6432 30010 6488
rect 30066 6432 30666 6488
rect 30005 6430 30666 6432
rect 30005 6427 30071 6430
rect 30465 6354 30531 6357
rect 28950 6352 30531 6354
rect 28950 6296 30470 6352
rect 30526 6296 30531 6352
rect 28950 6294 30531 6296
rect 30606 6354 30666 6430
rect 32673 6488 35959 6490
rect 32673 6432 32678 6488
rect 32734 6432 35898 6488
rect 35954 6432 35959 6488
rect 32673 6430 35959 6432
rect 32673 6427 32739 6430
rect 35893 6427 35959 6430
rect 36169 6354 36235 6357
rect 30606 6352 36235 6354
rect 30606 6296 36174 6352
rect 36230 6296 36235 6352
rect 30606 6294 36235 6296
rect 30465 6291 30531 6294
rect 36169 6291 36235 6294
rect 32581 6218 32647 6221
rect 35249 6218 35315 6221
rect 9860 6216 12591 6218
rect 9860 6160 12530 6216
rect 12586 6160 12591 6216
rect 9860 6158 12591 6160
rect 2681 5674 2747 5677
rect 3558 5674 3618 6158
rect 9581 6155 9647 6158
rect 12525 6155 12591 6158
rect 15104 6158 19350 6218
rect 22050 6216 32647 6218
rect 22050 6160 32586 6216
rect 32642 6160 32647 6216
rect 22050 6158 32647 6160
rect 13169 6082 13235 6085
rect 6134 6080 13235 6082
rect 6134 6024 13174 6080
rect 13230 6024 13235 6080
rect 6134 6022 13235 6024
rect 5707 6016 6023 6017
rect 5707 5952 5713 6016
rect 5777 5952 5793 6016
rect 5857 5952 5873 6016
rect 5937 5952 5953 6016
rect 6017 5952 6023 6016
rect 5707 5951 6023 5952
rect 4337 5810 4403 5813
rect 6134 5810 6194 6022
rect 13169 6019 13235 6022
rect 11605 5946 11671 5949
rect 14917 5946 14983 5949
rect 15104 5946 15164 6158
rect 15745 6082 15811 6085
rect 17585 6082 17651 6085
rect 15745 6080 17651 6082
rect 15745 6024 15750 6080
rect 15806 6024 17590 6080
rect 17646 6024 17651 6080
rect 15745 6022 17651 6024
rect 19290 6082 19350 6158
rect 32581 6155 32647 6158
rect 34148 6216 35315 6218
rect 34148 6160 35254 6216
rect 35310 6160 35315 6216
rect 34148 6158 35315 6160
rect 20805 6082 20871 6085
rect 22461 6082 22527 6085
rect 19290 6080 22527 6082
rect 19290 6024 20810 6080
rect 20866 6024 22466 6080
rect 22522 6024 22527 6080
rect 19290 6022 22527 6024
rect 15745 6019 15811 6022
rect 17585 6019 17651 6022
rect 20805 6019 20871 6022
rect 22461 6019 22527 6022
rect 25814 6020 25820 6084
rect 25884 6082 25890 6084
rect 34148 6082 34208 6158
rect 35249 6155 35315 6158
rect 25884 6022 34208 6082
rect 25884 6020 25890 6022
rect 15229 6016 15545 6017
rect 15229 5952 15235 6016
rect 15299 5952 15315 6016
rect 15379 5952 15395 6016
rect 15459 5952 15475 6016
rect 15539 5952 15545 6016
rect 15229 5951 15545 5952
rect 24751 6016 25067 6017
rect 24751 5952 24757 6016
rect 24821 5952 24837 6016
rect 24901 5952 24917 6016
rect 24981 5952 24997 6016
rect 25061 5952 25067 6016
rect 24751 5951 25067 5952
rect 34273 6016 34589 6017
rect 34273 5952 34279 6016
rect 34343 5952 34359 6016
rect 34423 5952 34439 6016
rect 34503 5952 34519 6016
rect 34583 5952 34589 6016
rect 34273 5951 34589 5952
rect 11605 5944 15164 5946
rect 11605 5888 11610 5944
rect 11666 5888 14922 5944
rect 14978 5888 15164 5944
rect 11605 5886 15164 5888
rect 15745 5946 15811 5949
rect 16205 5946 16271 5949
rect 20253 5946 20319 5949
rect 15745 5944 20319 5946
rect 15745 5888 15750 5944
rect 15806 5888 16210 5944
rect 16266 5888 20258 5944
rect 20314 5888 20319 5944
rect 15745 5886 20319 5888
rect 11605 5883 11671 5886
rect 14917 5883 14983 5886
rect 15745 5883 15811 5886
rect 16205 5883 16271 5886
rect 20253 5883 20319 5886
rect 21909 5946 21975 5949
rect 22093 5946 22159 5949
rect 25589 5948 25655 5949
rect 25589 5946 25636 5948
rect 21909 5944 22159 5946
rect 21909 5888 21914 5944
rect 21970 5888 22098 5944
rect 22154 5888 22159 5944
rect 21909 5886 22159 5888
rect 25544 5944 25636 5946
rect 25544 5888 25594 5944
rect 25544 5886 25636 5888
rect 21909 5883 21975 5886
rect 22093 5883 22159 5886
rect 25589 5884 25636 5886
rect 25700 5884 25706 5948
rect 26182 5884 26188 5948
rect 26252 5946 26258 5948
rect 26417 5946 26483 5949
rect 26252 5944 26483 5946
rect 26252 5888 26422 5944
rect 26478 5888 26483 5944
rect 26252 5886 26483 5888
rect 26252 5884 26258 5886
rect 25589 5883 25655 5884
rect 26417 5883 26483 5886
rect 27797 5946 27863 5949
rect 28533 5946 28599 5949
rect 27797 5944 28599 5946
rect 27797 5888 27802 5944
rect 27858 5888 28538 5944
rect 28594 5888 28599 5944
rect 27797 5886 28599 5888
rect 27797 5883 27863 5886
rect 28533 5883 28599 5886
rect 30414 5884 30420 5948
rect 30484 5946 30490 5948
rect 33961 5946 34027 5949
rect 30484 5944 34027 5946
rect 30484 5888 33966 5944
rect 34022 5888 34027 5944
rect 30484 5886 34027 5888
rect 30484 5884 30490 5886
rect 33961 5883 34027 5886
rect 4337 5808 6194 5810
rect 4337 5752 4342 5808
rect 4398 5752 6194 5808
rect 4337 5750 6194 5752
rect 10225 5810 10291 5813
rect 13261 5810 13327 5813
rect 15193 5810 15259 5813
rect 10225 5808 13327 5810
rect 10225 5752 10230 5808
rect 10286 5752 13266 5808
rect 13322 5752 13327 5808
rect 10225 5750 13327 5752
rect 4337 5747 4403 5750
rect 10225 5747 10291 5750
rect 13261 5747 13327 5750
rect 14046 5808 15259 5810
rect 14046 5752 15198 5808
rect 15254 5752 15259 5808
rect 14046 5750 15259 5752
rect 2681 5672 3618 5674
rect 2681 5616 2686 5672
rect 2742 5616 3618 5672
rect 2681 5614 3618 5616
rect 3693 5674 3759 5677
rect 9673 5676 9739 5677
rect 8886 5674 8892 5676
rect 3693 5672 8892 5674
rect 3693 5616 3698 5672
rect 3754 5616 8892 5672
rect 3693 5614 8892 5616
rect 2681 5611 2747 5614
rect 3693 5611 3759 5614
rect 8886 5612 8892 5614
rect 8956 5612 8962 5676
rect 9622 5612 9628 5676
rect 9692 5674 9739 5676
rect 9692 5672 9784 5674
rect 9734 5616 9784 5672
rect 9692 5614 9784 5616
rect 9692 5612 9739 5614
rect 11094 5612 11100 5676
rect 11164 5674 11170 5676
rect 14046 5674 14106 5750
rect 15193 5747 15259 5750
rect 19609 5810 19675 5813
rect 28257 5810 28323 5813
rect 19609 5808 28323 5810
rect 19609 5752 19614 5808
rect 19670 5752 28262 5808
rect 28318 5752 28323 5808
rect 19609 5750 28323 5752
rect 19609 5747 19675 5750
rect 28257 5747 28323 5750
rect 28625 5810 28691 5813
rect 28625 5808 29332 5810
rect 28625 5752 28630 5808
rect 28686 5752 29332 5808
rect 28625 5750 29332 5752
rect 28625 5747 28691 5750
rect 11164 5614 14106 5674
rect 14733 5674 14799 5677
rect 24761 5674 24827 5677
rect 28441 5674 28507 5677
rect 14733 5672 21144 5674
rect 14733 5616 14738 5672
rect 14794 5616 21144 5672
rect 14733 5614 21144 5616
rect 11164 5612 11170 5614
rect 9673 5611 9739 5612
rect 14733 5611 14799 5614
rect 0 5538 800 5568
rect 21084 5541 21144 5614
rect 24761 5672 28507 5674
rect 24761 5616 24766 5672
rect 24822 5616 28446 5672
rect 28502 5616 28507 5672
rect 24761 5614 28507 5616
rect 24761 5611 24827 5614
rect 28441 5611 28507 5614
rect 29272 5541 29332 5750
rect 30373 5674 30439 5677
rect 33317 5674 33383 5677
rect 33593 5674 33659 5677
rect 30373 5672 33659 5674
rect 30373 5616 30378 5672
rect 30434 5616 33322 5672
rect 33378 5616 33598 5672
rect 33654 5616 33659 5672
rect 30373 5614 33659 5616
rect 30373 5611 30439 5614
rect 33317 5611 33383 5614
rect 33593 5611 33659 5614
rect 1025 5538 1091 5541
rect 0 5536 1091 5538
rect 0 5480 1030 5536
rect 1086 5480 1091 5536
rect 0 5478 1091 5480
rect 0 5448 800 5478
rect 1025 5475 1091 5478
rect 4521 5538 4587 5541
rect 9121 5538 9187 5541
rect 4521 5536 9187 5538
rect 4521 5480 4526 5536
rect 4582 5480 9126 5536
rect 9182 5480 9187 5536
rect 4521 5478 9187 5480
rect 4521 5475 4587 5478
rect 9121 5475 9187 5478
rect 14273 5538 14339 5541
rect 15377 5538 15443 5541
rect 14273 5536 15443 5538
rect 14273 5480 14278 5536
rect 14334 5480 15382 5536
rect 15438 5480 15443 5536
rect 14273 5478 15443 5480
rect 14273 5475 14339 5478
rect 15377 5475 15443 5478
rect 15561 5538 15627 5541
rect 16665 5540 16731 5541
rect 15878 5538 15884 5540
rect 15561 5536 15884 5538
rect 15561 5480 15566 5536
rect 15622 5480 15884 5536
rect 15561 5478 15884 5480
rect 15561 5475 15627 5478
rect 15878 5476 15884 5478
rect 15948 5476 15954 5540
rect 16614 5538 16620 5540
rect 16574 5478 16620 5538
rect 16684 5536 16731 5540
rect 16726 5480 16731 5536
rect 16614 5476 16620 5478
rect 16684 5476 16731 5480
rect 16665 5475 16731 5476
rect 21081 5538 21147 5541
rect 27613 5538 27679 5541
rect 21081 5536 27679 5538
rect 21081 5480 21086 5536
rect 21142 5480 27618 5536
rect 27674 5480 27679 5536
rect 21081 5478 27679 5480
rect 21081 5475 21147 5478
rect 27613 5475 27679 5478
rect 27797 5538 27863 5541
rect 27797 5536 29010 5538
rect 27797 5480 27802 5536
rect 27858 5480 29010 5536
rect 27797 5478 29010 5480
rect 27797 5475 27863 5478
rect 10468 5472 10784 5473
rect 10468 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10784 5472
rect 10468 5407 10784 5408
rect 19990 5472 20306 5473
rect 19990 5408 19996 5472
rect 20060 5408 20076 5472
rect 20140 5408 20156 5472
rect 20220 5408 20236 5472
rect 20300 5408 20306 5472
rect 19990 5407 20306 5408
rect 5993 5402 6059 5405
rect 6310 5402 6316 5404
rect 5993 5400 6316 5402
rect 5993 5344 5998 5400
rect 6054 5344 6316 5400
rect 5993 5342 6316 5344
rect 5993 5339 6059 5342
rect 6310 5340 6316 5342
rect 6380 5340 6386 5404
rect 13302 5340 13308 5404
rect 13372 5402 13378 5404
rect 22369 5402 22435 5405
rect 23013 5402 23079 5405
rect 13372 5342 16314 5402
rect 13372 5340 13378 5342
rect 2814 5204 2820 5268
rect 2884 5266 2890 5268
rect 15285 5266 15351 5269
rect 2884 5264 15351 5266
rect 2884 5208 15290 5264
rect 15346 5208 15351 5264
rect 2884 5206 15351 5208
rect 2884 5204 2890 5206
rect 15285 5203 15351 5206
rect 15469 5266 15535 5269
rect 16113 5266 16179 5269
rect 15469 5264 16179 5266
rect 15469 5208 15474 5264
rect 15530 5208 16118 5264
rect 16174 5208 16179 5264
rect 15469 5206 16179 5208
rect 16254 5266 16314 5342
rect 22369 5400 23079 5402
rect 22369 5344 22374 5400
rect 22430 5344 23018 5400
rect 23074 5344 23079 5400
rect 22369 5342 23079 5344
rect 22369 5339 22435 5342
rect 23013 5339 23079 5342
rect 22461 5266 22527 5269
rect 25497 5266 25563 5269
rect 16254 5264 25563 5266
rect 16254 5208 22466 5264
rect 22522 5208 25502 5264
rect 25558 5208 25563 5264
rect 16254 5206 25563 5208
rect 15469 5203 15535 5206
rect 16113 5203 16179 5206
rect 22461 5203 22527 5206
rect 25497 5203 25563 5206
rect 27429 5266 27495 5269
rect 28206 5266 28212 5268
rect 27429 5264 28212 5266
rect 27429 5208 27434 5264
rect 27490 5208 28212 5264
rect 27429 5206 28212 5208
rect 27429 5203 27495 5206
rect 28206 5204 28212 5206
rect 28276 5266 28282 5268
rect 28441 5266 28507 5269
rect 28276 5264 28507 5266
rect 28276 5208 28446 5264
rect 28502 5208 28507 5264
rect 28276 5206 28507 5208
rect 28950 5266 29010 5478
rect 29269 5536 29335 5541
rect 29269 5480 29274 5536
rect 29330 5480 29335 5536
rect 29269 5475 29335 5480
rect 33593 5538 33659 5541
rect 33726 5538 33732 5540
rect 33593 5536 33732 5538
rect 33593 5480 33598 5536
rect 33654 5480 33732 5536
rect 33593 5478 33732 5480
rect 33593 5475 33659 5478
rect 33726 5476 33732 5478
rect 33796 5476 33802 5540
rect 29512 5472 29828 5473
rect 29512 5408 29518 5472
rect 29582 5408 29598 5472
rect 29662 5408 29678 5472
rect 29742 5408 29758 5472
rect 29822 5408 29828 5472
rect 29512 5407 29828 5408
rect 39034 5472 39350 5473
rect 39034 5408 39040 5472
rect 39104 5408 39120 5472
rect 39184 5408 39200 5472
rect 39264 5408 39280 5472
rect 39344 5408 39350 5472
rect 39566 5448 40366 5568
rect 39034 5407 39350 5408
rect 29913 5402 29979 5405
rect 31017 5402 31083 5405
rect 29913 5400 31083 5402
rect 29913 5344 29918 5400
rect 29974 5344 31022 5400
rect 31078 5344 31083 5400
rect 29913 5342 31083 5344
rect 29913 5339 29979 5342
rect 31017 5339 31083 5342
rect 30465 5266 30531 5269
rect 28950 5264 30531 5266
rect 28950 5208 30470 5264
rect 30526 5208 30531 5264
rect 28950 5206 30531 5208
rect 28276 5204 28282 5206
rect 28441 5203 28507 5206
rect 30465 5203 30531 5206
rect 31109 5266 31175 5269
rect 36813 5266 36879 5269
rect 31109 5264 36879 5266
rect 31109 5208 31114 5264
rect 31170 5208 36818 5264
rect 36874 5208 36879 5264
rect 31109 5206 36879 5208
rect 31109 5203 31175 5206
rect 36813 5203 36879 5206
rect 5349 5130 5415 5133
rect 14825 5130 14891 5133
rect 5349 5128 14891 5130
rect 5349 5072 5354 5128
rect 5410 5072 14830 5128
rect 14886 5072 14891 5128
rect 5349 5070 14891 5072
rect 5349 5067 5415 5070
rect 14825 5067 14891 5070
rect 15009 5130 15075 5133
rect 20989 5130 21055 5133
rect 15009 5128 21055 5130
rect 15009 5072 15014 5128
rect 15070 5072 20994 5128
rect 21050 5072 21055 5128
rect 15009 5070 21055 5072
rect 15009 5067 15075 5070
rect 20989 5067 21055 5070
rect 26785 5130 26851 5133
rect 36905 5130 36971 5133
rect 26785 5128 36971 5130
rect 26785 5072 26790 5128
rect 26846 5072 36910 5128
rect 36966 5072 36971 5128
rect 26785 5070 36971 5072
rect 26785 5067 26851 5070
rect 36905 5067 36971 5070
rect 7598 4932 7604 4996
rect 7668 4994 7674 4996
rect 14365 4994 14431 4997
rect 7668 4992 14431 4994
rect 7668 4936 14370 4992
rect 14426 4936 14431 4992
rect 7668 4934 14431 4936
rect 7668 4932 7674 4934
rect 14365 4931 14431 4934
rect 19517 4994 19583 4997
rect 23841 4994 23907 4997
rect 19517 4992 23907 4994
rect 19517 4936 19522 4992
rect 19578 4936 23846 4992
rect 23902 4936 23907 4992
rect 19517 4934 23907 4936
rect 19517 4931 19583 4934
rect 23841 4931 23907 4934
rect 25773 4994 25839 4997
rect 32397 4994 32463 4997
rect 25773 4992 32463 4994
rect 25773 4936 25778 4992
rect 25834 4936 32402 4992
rect 32458 4936 32463 4992
rect 25773 4934 32463 4936
rect 25773 4931 25839 4934
rect 32397 4931 32463 4934
rect 5707 4928 6023 4929
rect 5707 4864 5713 4928
rect 5777 4864 5793 4928
rect 5857 4864 5873 4928
rect 5937 4864 5953 4928
rect 6017 4864 6023 4928
rect 5707 4863 6023 4864
rect 15229 4928 15545 4929
rect 15229 4864 15235 4928
rect 15299 4864 15315 4928
rect 15379 4864 15395 4928
rect 15459 4864 15475 4928
rect 15539 4864 15545 4928
rect 15229 4863 15545 4864
rect 24751 4928 25067 4929
rect 24751 4864 24757 4928
rect 24821 4864 24837 4928
rect 24901 4864 24917 4928
rect 24981 4864 24997 4928
rect 25061 4864 25067 4928
rect 24751 4863 25067 4864
rect 34273 4928 34589 4929
rect 34273 4864 34279 4928
rect 34343 4864 34359 4928
rect 34423 4864 34439 4928
rect 34503 4864 34519 4928
rect 34583 4864 34589 4928
rect 34273 4863 34589 4864
rect 6085 4858 6151 4861
rect 6637 4858 6703 4861
rect 8569 4858 8635 4861
rect 6085 4856 8635 4858
rect 6085 4800 6090 4856
rect 6146 4800 6642 4856
rect 6698 4800 8574 4856
rect 8630 4800 8635 4856
rect 6085 4798 8635 4800
rect 6085 4795 6151 4798
rect 6637 4795 6703 4798
rect 8569 4795 8635 4798
rect 10869 4858 10935 4861
rect 12249 4858 12315 4861
rect 13353 4860 13419 4861
rect 10869 4856 12315 4858
rect 10869 4800 10874 4856
rect 10930 4800 12254 4856
rect 12310 4800 12315 4856
rect 10869 4798 12315 4800
rect 10869 4795 10935 4798
rect 12249 4795 12315 4798
rect 13302 4796 13308 4860
rect 13372 4858 13419 4860
rect 28809 4858 28875 4861
rect 13372 4856 13464 4858
rect 13414 4800 13464 4856
rect 13372 4798 13464 4800
rect 26190 4856 28875 4858
rect 26190 4800 28814 4856
rect 28870 4800 28875 4856
rect 26190 4798 28875 4800
rect 13372 4796 13419 4798
rect 13353 4795 13419 4796
rect 5809 4722 5875 4725
rect 16297 4722 16363 4725
rect 5809 4720 16363 4722
rect 5809 4664 5814 4720
rect 5870 4664 16302 4720
rect 16358 4664 16363 4720
rect 5809 4662 16363 4664
rect 5809 4659 5875 4662
rect 16297 4659 16363 4662
rect 7465 4586 7531 4589
rect 14549 4586 14615 4589
rect 26190 4586 26250 4798
rect 28809 4795 28875 4798
rect 30741 4858 30807 4861
rect 33777 4858 33843 4861
rect 30741 4856 33843 4858
rect 30741 4800 30746 4856
rect 30802 4800 33782 4856
rect 33838 4800 33843 4856
rect 30741 4798 33843 4800
rect 30741 4795 30807 4798
rect 33777 4795 33843 4798
rect 26325 4722 26391 4725
rect 35433 4722 35499 4725
rect 26325 4720 35499 4722
rect 26325 4664 26330 4720
rect 26386 4664 35438 4720
rect 35494 4664 35499 4720
rect 26325 4662 35499 4664
rect 26325 4659 26391 4662
rect 35433 4659 35499 4662
rect 31661 4586 31727 4589
rect 7465 4584 12450 4586
rect 7465 4528 7470 4584
rect 7526 4528 12450 4584
rect 7465 4526 12450 4528
rect 7465 4523 7531 4526
rect 12390 4450 12450 4526
rect 14549 4584 26250 4586
rect 14549 4528 14554 4584
rect 14610 4528 26250 4584
rect 14549 4526 26250 4528
rect 27294 4584 31727 4586
rect 27294 4528 31666 4584
rect 31722 4528 31727 4584
rect 27294 4526 31727 4528
rect 14549 4523 14615 4526
rect 18781 4450 18847 4453
rect 12390 4448 18847 4450
rect 12390 4392 18786 4448
rect 18842 4392 18847 4448
rect 12390 4390 18847 4392
rect 18781 4387 18847 4390
rect 19333 4450 19399 4453
rect 19517 4450 19583 4453
rect 19333 4448 19583 4450
rect 19333 4392 19338 4448
rect 19394 4392 19522 4448
rect 19578 4392 19583 4448
rect 19333 4390 19583 4392
rect 19333 4387 19399 4390
rect 19517 4387 19583 4390
rect 26325 4450 26391 4453
rect 27102 4450 27108 4452
rect 26325 4448 27108 4450
rect 26325 4392 26330 4448
rect 26386 4392 27108 4448
rect 26325 4390 27108 4392
rect 26325 4387 26391 4390
rect 27102 4388 27108 4390
rect 27172 4388 27178 4452
rect 10468 4384 10784 4385
rect 10468 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10784 4384
rect 10468 4319 10784 4320
rect 19990 4384 20306 4385
rect 19990 4320 19996 4384
rect 20060 4320 20076 4384
rect 20140 4320 20156 4384
rect 20220 4320 20236 4384
rect 20300 4320 20306 4384
rect 19990 4319 20306 4320
rect 2773 4314 2839 4317
rect 10317 4314 10383 4317
rect 2773 4312 10383 4314
rect 2773 4256 2778 4312
rect 2834 4256 10322 4312
rect 10378 4256 10383 4312
rect 2773 4254 10383 4256
rect 2773 4251 2839 4254
rect 10317 4251 10383 4254
rect 15561 4314 15627 4317
rect 18321 4314 18387 4317
rect 19517 4314 19583 4317
rect 15561 4312 19583 4314
rect 15561 4256 15566 4312
rect 15622 4256 18326 4312
rect 18382 4256 19522 4312
rect 19578 4256 19583 4312
rect 15561 4254 19583 4256
rect 15561 4251 15627 4254
rect 18321 4251 18387 4254
rect 19517 4251 19583 4254
rect 4521 4178 4587 4181
rect 5206 4178 5212 4180
rect 4521 4176 5212 4178
rect 4521 4120 4526 4176
rect 4582 4120 5212 4176
rect 4521 4118 5212 4120
rect 4521 4115 4587 4118
rect 5206 4116 5212 4118
rect 5276 4116 5282 4180
rect 10133 4178 10199 4181
rect 10685 4178 10751 4181
rect 10133 4176 10751 4178
rect 10133 4120 10138 4176
rect 10194 4120 10690 4176
rect 10746 4120 10751 4176
rect 10133 4118 10751 4120
rect 10133 4115 10199 4118
rect 10685 4115 10751 4118
rect 13169 4178 13235 4181
rect 16297 4178 16363 4181
rect 27294 4178 27354 4526
rect 31661 4523 31727 4526
rect 29512 4384 29828 4385
rect 29512 4320 29518 4384
rect 29582 4320 29598 4384
rect 29662 4320 29678 4384
rect 29742 4320 29758 4384
rect 29822 4320 29828 4384
rect 29512 4319 29828 4320
rect 39034 4384 39350 4385
rect 39034 4320 39040 4384
rect 39104 4320 39120 4384
rect 39184 4320 39200 4384
rect 39264 4320 39280 4384
rect 39344 4320 39350 4384
rect 39034 4319 39350 4320
rect 37641 4178 37707 4181
rect 13169 4176 27354 4178
rect 13169 4120 13174 4176
rect 13230 4120 16302 4176
rect 16358 4120 27354 4176
rect 13169 4118 27354 4120
rect 28950 4176 37707 4178
rect 28950 4120 37646 4176
rect 37702 4120 37707 4176
rect 28950 4118 37707 4120
rect 13169 4115 13235 4118
rect 16297 4115 16363 4118
rect 3969 4042 4035 4045
rect 5717 4042 5783 4045
rect 3969 4040 5783 4042
rect 3969 3984 3974 4040
rect 4030 3984 5722 4040
rect 5778 3984 5783 4040
rect 3969 3982 5783 3984
rect 3969 3979 4035 3982
rect 5717 3979 5783 3982
rect 5901 4042 5967 4045
rect 7925 4042 7991 4045
rect 12249 4044 12315 4045
rect 17953 4044 18019 4045
rect 12198 4042 12204 4044
rect 5901 4040 7991 4042
rect 5901 3984 5906 4040
rect 5962 3984 7930 4040
rect 7986 3984 7991 4040
rect 5901 3982 7991 3984
rect 12158 3982 12204 4042
rect 12268 4040 12315 4044
rect 17902 4042 17908 4044
rect 12310 3984 12315 4040
rect 5901 3979 5967 3982
rect 5707 3840 6023 3841
rect 5707 3776 5713 3840
rect 5777 3776 5793 3840
rect 5857 3776 5873 3840
rect 5937 3776 5953 3840
rect 6017 3776 6023 3840
rect 5707 3775 6023 3776
rect 1853 3634 1919 3637
rect 3182 3634 3188 3636
rect 1853 3632 3188 3634
rect 1853 3576 1858 3632
rect 1914 3576 3188 3632
rect 1853 3574 3188 3576
rect 1853 3571 1919 3574
rect 3182 3572 3188 3574
rect 3252 3572 3258 3636
rect 3509 3634 3575 3637
rect 4797 3634 4863 3637
rect 6134 3634 6194 3982
rect 7925 3979 7991 3982
rect 12198 3980 12204 3982
rect 12268 3980 12315 3984
rect 12249 3979 12315 3980
rect 12390 3982 17050 4042
rect 17862 3982 17908 4042
rect 17972 4040 18019 4044
rect 18014 3984 18019 4040
rect 12014 3844 12020 3908
rect 12084 3906 12090 3908
rect 12390 3906 12450 3982
rect 12084 3846 12450 3906
rect 16990 3906 17050 3982
rect 17902 3980 17908 3982
rect 17972 3980 18019 3984
rect 17953 3979 18019 3980
rect 18229 4044 18295 4045
rect 18229 4040 18276 4044
rect 18340 4042 18346 4044
rect 21357 4042 21423 4045
rect 26049 4042 26115 4045
rect 28950 4042 29010 4118
rect 37641 4115 37707 4118
rect 18229 3984 18234 4040
rect 18229 3980 18276 3984
rect 18340 3982 18386 4042
rect 21357 4040 25192 4042
rect 21357 3984 21362 4040
rect 21418 3984 25192 4040
rect 21357 3982 25192 3984
rect 18340 3980 18346 3982
rect 18229 3979 18295 3980
rect 21357 3979 21423 3982
rect 25132 3909 25192 3982
rect 26049 4040 29010 4042
rect 26049 3984 26054 4040
rect 26110 3984 29010 4040
rect 26049 3982 29010 3984
rect 30005 4044 30071 4045
rect 30005 4040 30052 4044
rect 30116 4042 30122 4044
rect 31385 4042 31451 4045
rect 36261 4042 36327 4045
rect 30005 3984 30010 4040
rect 26049 3979 26115 3982
rect 30005 3980 30052 3984
rect 30116 3982 30162 4042
rect 31385 4040 36327 4042
rect 31385 3984 31390 4040
rect 31446 3984 36266 4040
rect 36322 3984 36327 4040
rect 31385 3982 36327 3984
rect 30116 3980 30122 3982
rect 30005 3979 30071 3980
rect 31385 3979 31451 3982
rect 36261 3979 36327 3982
rect 21081 3906 21147 3909
rect 16990 3904 21147 3906
rect 16990 3848 21086 3904
rect 21142 3848 21147 3904
rect 16990 3846 21147 3848
rect 12084 3844 12090 3846
rect 21081 3843 21147 3846
rect 25129 3906 25195 3909
rect 25957 3906 26023 3909
rect 31569 3906 31635 3909
rect 32397 3906 32463 3909
rect 32673 3908 32739 3909
rect 32622 3906 32628 3908
rect 25129 3904 32463 3906
rect 25129 3848 25134 3904
rect 25190 3848 25962 3904
rect 26018 3848 31574 3904
rect 31630 3848 32402 3904
rect 32458 3848 32463 3904
rect 25129 3846 32463 3848
rect 32582 3846 32628 3906
rect 32692 3904 32739 3908
rect 32734 3848 32739 3904
rect 25129 3843 25195 3846
rect 25957 3843 26023 3846
rect 31569 3843 31635 3846
rect 32397 3843 32463 3846
rect 32622 3844 32628 3846
rect 32692 3844 32739 3848
rect 32673 3843 32739 3844
rect 15229 3840 15545 3841
rect 15229 3776 15235 3840
rect 15299 3776 15315 3840
rect 15379 3776 15395 3840
rect 15459 3776 15475 3840
rect 15539 3776 15545 3840
rect 15229 3775 15545 3776
rect 24751 3840 25067 3841
rect 24751 3776 24757 3840
rect 24821 3776 24837 3840
rect 24901 3776 24917 3840
rect 24981 3776 24997 3840
rect 25061 3776 25067 3840
rect 24751 3775 25067 3776
rect 34273 3840 34589 3841
rect 34273 3776 34279 3840
rect 34343 3776 34359 3840
rect 34423 3776 34439 3840
rect 34503 3776 34519 3840
rect 34583 3776 34589 3840
rect 34273 3775 34589 3776
rect 27429 3770 27495 3773
rect 25132 3768 27495 3770
rect 25132 3712 27434 3768
rect 27490 3712 27495 3768
rect 25132 3710 27495 3712
rect 3509 3632 6194 3634
rect 3509 3576 3514 3632
rect 3570 3576 4802 3632
rect 4858 3576 6194 3632
rect 3509 3574 6194 3576
rect 11237 3634 11303 3637
rect 25132 3634 25192 3710
rect 27429 3707 27495 3710
rect 36629 3634 36695 3637
rect 11237 3632 25192 3634
rect 11237 3576 11242 3632
rect 11298 3576 25192 3632
rect 11237 3574 25192 3576
rect 26006 3632 36695 3634
rect 26006 3576 36634 3632
rect 36690 3576 36695 3632
rect 26006 3574 36695 3576
rect 3509 3571 3575 3574
rect 4797 3571 4863 3574
rect 11237 3571 11303 3574
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 5993 3498 6059 3501
rect 13445 3498 13511 3501
rect 17033 3498 17099 3501
rect 26006 3498 26066 3574
rect 36629 3571 36695 3574
rect 5993 3496 12450 3498
rect 5993 3440 5998 3496
rect 6054 3440 12450 3496
rect 5993 3438 12450 3440
rect 5993 3435 6059 3438
rect 5717 3362 5783 3365
rect 7833 3362 7899 3365
rect 5717 3360 7899 3362
rect 5717 3304 5722 3360
rect 5778 3304 7838 3360
rect 7894 3304 7899 3360
rect 5717 3302 7899 3304
rect 12390 3362 12450 3438
rect 13445 3496 17099 3498
rect 13445 3440 13450 3496
rect 13506 3440 17038 3496
rect 17094 3440 17099 3496
rect 13445 3438 17099 3440
rect 13445 3435 13511 3438
rect 17033 3435 17099 3438
rect 17174 3438 26066 3498
rect 26141 3498 26207 3501
rect 38653 3498 38719 3501
rect 39566 3498 40366 3528
rect 26141 3496 31770 3498
rect 26141 3440 26146 3496
rect 26202 3440 31770 3496
rect 26141 3438 31770 3440
rect 17174 3362 17234 3438
rect 26141 3435 26207 3438
rect 12390 3302 17234 3362
rect 23381 3362 23447 3365
rect 28942 3362 28948 3364
rect 23381 3360 28948 3362
rect 23381 3304 23386 3360
rect 23442 3304 28948 3360
rect 23381 3302 28948 3304
rect 5717 3299 5783 3302
rect 7833 3299 7899 3302
rect 23381 3299 23447 3302
rect 28942 3300 28948 3302
rect 29012 3300 29018 3364
rect 31710 3362 31770 3438
rect 38653 3496 40366 3498
rect 38653 3440 38658 3496
rect 38714 3440 40366 3496
rect 38653 3438 40366 3440
rect 38653 3435 38719 3438
rect 39566 3408 40366 3438
rect 34646 3362 34652 3364
rect 31710 3302 34652 3362
rect 34646 3300 34652 3302
rect 34716 3300 34722 3364
rect 10468 3296 10784 3297
rect 10468 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10784 3296
rect 10468 3231 10784 3232
rect 19990 3296 20306 3297
rect 19990 3232 19996 3296
rect 20060 3232 20076 3296
rect 20140 3232 20156 3296
rect 20220 3232 20236 3296
rect 20300 3232 20306 3296
rect 19990 3231 20306 3232
rect 29512 3296 29828 3297
rect 29512 3232 29518 3296
rect 29582 3232 29598 3296
rect 29662 3232 29678 3296
rect 29742 3232 29758 3296
rect 29822 3232 29828 3296
rect 29512 3231 29828 3232
rect 39034 3296 39350 3297
rect 39034 3232 39040 3296
rect 39104 3232 39120 3296
rect 39184 3232 39200 3296
rect 39264 3232 39280 3296
rect 39344 3232 39350 3296
rect 39034 3231 39350 3232
rect 1853 3226 1919 3229
rect 7281 3226 7347 3229
rect 1853 3224 7347 3226
rect 1853 3168 1858 3224
rect 1914 3168 7286 3224
rect 7342 3168 7347 3224
rect 1853 3166 7347 3168
rect 1853 3163 1919 3166
rect 7281 3163 7347 3166
rect 11053 3226 11119 3229
rect 13445 3226 13511 3229
rect 11053 3224 13511 3226
rect 11053 3168 11058 3224
rect 11114 3168 13450 3224
rect 13506 3168 13511 3224
rect 11053 3166 13511 3168
rect 11053 3163 11119 3166
rect 13445 3163 13511 3166
rect 13905 3226 13971 3229
rect 26601 3226 26667 3229
rect 26734 3226 26740 3228
rect 13905 3224 14290 3226
rect 13905 3168 13910 3224
rect 13966 3168 14290 3224
rect 13905 3166 14290 3168
rect 13905 3163 13971 3166
rect 5717 3090 5783 3093
rect 14089 3092 14155 3093
rect 14038 3090 14044 3092
rect 5717 3088 14044 3090
rect 14108 3088 14155 3092
rect 5717 3032 5722 3088
rect 5778 3032 14044 3088
rect 14150 3032 14155 3088
rect 5717 3030 14044 3032
rect 5717 3027 5783 3030
rect 14038 3028 14044 3030
rect 14108 3028 14155 3032
rect 14230 3090 14290 3166
rect 26601 3224 26740 3226
rect 26601 3168 26606 3224
rect 26662 3168 26740 3224
rect 26601 3166 26740 3168
rect 26601 3163 26667 3166
rect 26734 3164 26740 3166
rect 26804 3226 26810 3228
rect 27521 3226 27587 3229
rect 26804 3224 27587 3226
rect 26804 3168 27526 3224
rect 27582 3168 27587 3224
rect 26804 3166 27587 3168
rect 26804 3164 26810 3166
rect 27521 3163 27587 3166
rect 21449 3090 21515 3093
rect 33409 3090 33475 3093
rect 14230 3030 21098 3090
rect 14089 3027 14155 3028
rect 4797 2954 4863 2957
rect 6637 2954 6703 2957
rect 20897 2954 20963 2957
rect 4797 2952 6194 2954
rect 4797 2896 4802 2952
rect 4858 2896 6194 2952
rect 4797 2894 6194 2896
rect 4797 2891 4863 2894
rect 6134 2818 6194 2894
rect 6637 2952 20963 2954
rect 6637 2896 6642 2952
rect 6698 2896 20902 2952
rect 20958 2896 20963 2952
rect 6637 2894 20963 2896
rect 21038 2954 21098 3030
rect 21449 3088 33475 3090
rect 21449 3032 21454 3088
rect 21510 3032 33414 3088
rect 33470 3032 33475 3088
rect 21449 3030 33475 3032
rect 21449 3027 21515 3030
rect 33409 3027 33475 3030
rect 36813 2954 36879 2957
rect 21038 2952 36879 2954
rect 21038 2896 36818 2952
rect 36874 2896 36879 2952
rect 21038 2894 36879 2896
rect 6637 2891 6703 2894
rect 20897 2891 20963 2894
rect 36813 2891 36879 2894
rect 6913 2818 6979 2821
rect 6134 2816 6979 2818
rect 6134 2760 6918 2816
rect 6974 2760 6979 2816
rect 6134 2758 6979 2760
rect 6913 2755 6979 2758
rect 17033 2818 17099 2821
rect 19425 2818 19491 2821
rect 21909 2818 21975 2821
rect 17033 2816 21975 2818
rect 17033 2760 17038 2816
rect 17094 2760 19430 2816
rect 19486 2760 21914 2816
rect 21970 2760 21975 2816
rect 17033 2758 21975 2760
rect 17033 2755 17099 2758
rect 19425 2755 19491 2758
rect 21909 2755 21975 2758
rect 27429 2818 27495 2821
rect 31753 2818 31819 2821
rect 34145 2818 34211 2821
rect 27429 2816 34211 2818
rect 27429 2760 27434 2816
rect 27490 2760 31758 2816
rect 31814 2760 34150 2816
rect 34206 2760 34211 2816
rect 27429 2758 34211 2760
rect 27429 2755 27495 2758
rect 31753 2755 31819 2758
rect 34145 2755 34211 2758
rect 5707 2752 6023 2753
rect 5707 2688 5713 2752
rect 5777 2688 5793 2752
rect 5857 2688 5873 2752
rect 5937 2688 5953 2752
rect 6017 2688 6023 2752
rect 5707 2687 6023 2688
rect 15229 2752 15545 2753
rect 15229 2688 15235 2752
rect 15299 2688 15315 2752
rect 15379 2688 15395 2752
rect 15459 2688 15475 2752
rect 15539 2688 15545 2752
rect 15229 2687 15545 2688
rect 24751 2752 25067 2753
rect 24751 2688 24757 2752
rect 24821 2688 24837 2752
rect 24901 2688 24917 2752
rect 24981 2688 24997 2752
rect 25061 2688 25067 2752
rect 24751 2687 25067 2688
rect 34273 2752 34589 2753
rect 34273 2688 34279 2752
rect 34343 2688 34359 2752
rect 34423 2688 34439 2752
rect 34503 2688 34519 2752
rect 34583 2688 34589 2752
rect 34273 2687 34589 2688
rect 17125 2684 17191 2685
rect 17125 2680 17172 2684
rect 17236 2682 17242 2684
rect 25129 2682 25195 2685
rect 33225 2684 33291 2685
rect 27654 2682 27660 2684
rect 17125 2624 17130 2680
rect 17125 2620 17172 2624
rect 17236 2622 17282 2682
rect 25129 2680 27660 2682
rect 25129 2624 25134 2680
rect 25190 2624 27660 2680
rect 25129 2622 27660 2624
rect 17236 2620 17242 2622
rect 17125 2619 17191 2620
rect 25129 2619 25195 2622
rect 27654 2620 27660 2622
rect 27724 2620 27730 2684
rect 33174 2682 33180 2684
rect 33134 2622 33180 2682
rect 33244 2680 33291 2684
rect 33286 2624 33291 2680
rect 33174 2620 33180 2622
rect 33244 2620 33291 2624
rect 33225 2619 33291 2620
rect 5390 2484 5396 2548
rect 5460 2546 5466 2548
rect 15193 2546 15259 2549
rect 18689 2546 18755 2549
rect 5460 2544 15259 2546
rect 5460 2488 15198 2544
rect 15254 2488 15259 2544
rect 5460 2486 15259 2488
rect 5460 2484 5466 2486
rect 15193 2483 15259 2486
rect 16530 2544 18755 2546
rect 16530 2488 18694 2544
rect 18750 2488 18755 2544
rect 16530 2486 18755 2488
rect 9765 2410 9831 2413
rect 16530 2410 16590 2486
rect 18689 2483 18755 2486
rect 23974 2484 23980 2548
rect 24044 2546 24050 2548
rect 25313 2546 25379 2549
rect 24044 2544 25379 2546
rect 24044 2488 25318 2544
rect 25374 2488 25379 2544
rect 24044 2486 25379 2488
rect 24044 2484 24050 2486
rect 25313 2483 25379 2486
rect 38469 2410 38535 2413
rect 9765 2408 16590 2410
rect 9765 2352 9770 2408
rect 9826 2352 16590 2408
rect 9765 2350 16590 2352
rect 19750 2408 38535 2410
rect 19750 2352 38474 2408
rect 38530 2352 38535 2408
rect 19750 2350 38535 2352
rect 9765 2347 9831 2350
rect 13813 2274 13879 2277
rect 19149 2274 19215 2277
rect 13813 2272 19215 2274
rect 13813 2216 13818 2272
rect 13874 2216 19154 2272
rect 19210 2216 19215 2272
rect 13813 2214 19215 2216
rect 13813 2211 13879 2214
rect 19149 2211 19215 2214
rect 10468 2208 10784 2209
rect 10468 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10784 2208
rect 10468 2143 10784 2144
rect 13629 2138 13695 2141
rect 19750 2138 19810 2350
rect 38469 2347 38535 2350
rect 19990 2208 20306 2209
rect 19990 2144 19996 2208
rect 20060 2144 20076 2208
rect 20140 2144 20156 2208
rect 20220 2144 20236 2208
rect 20300 2144 20306 2208
rect 19990 2143 20306 2144
rect 29512 2208 29828 2209
rect 29512 2144 29518 2208
rect 29582 2144 29598 2208
rect 29662 2144 29678 2208
rect 29742 2144 29758 2208
rect 29822 2144 29828 2208
rect 29512 2143 29828 2144
rect 39034 2208 39350 2209
rect 39034 2144 39040 2208
rect 39104 2144 39120 2208
rect 39184 2144 39200 2208
rect 39264 2144 39280 2208
rect 39344 2144 39350 2208
rect 39034 2143 39350 2144
rect 39566 2138 40366 2168
rect 13629 2136 19810 2138
rect 13629 2080 13634 2136
rect 13690 2080 19810 2136
rect 13629 2078 19810 2080
rect 39438 2078 40366 2138
rect 13629 2075 13695 2078
rect 7741 2002 7807 2005
rect 37273 2002 37339 2005
rect 7741 2000 37339 2002
rect 7741 1944 7746 2000
rect 7802 1944 37278 2000
rect 37334 1944 37339 2000
rect 7741 1942 37339 1944
rect 7741 1939 7807 1942
rect 37273 1939 37339 1942
rect 38653 2002 38719 2005
rect 39438 2002 39498 2078
rect 39566 2048 40366 2078
rect 38653 2000 39498 2002
rect 38653 1944 38658 2000
rect 38714 1944 39498 2000
rect 38653 1942 39498 1944
rect 38653 1939 38719 1942
rect 10174 1804 10180 1868
rect 10244 1866 10250 1868
rect 35893 1866 35959 1869
rect 10244 1864 35959 1866
rect 10244 1808 35898 1864
rect 35954 1808 35959 1864
rect 10244 1806 35959 1808
rect 10244 1804 10250 1806
rect 35893 1803 35959 1806
rect 13261 1730 13327 1733
rect 38193 1730 38259 1733
rect 13261 1728 38259 1730
rect 13261 1672 13266 1728
rect 13322 1672 38198 1728
rect 38254 1672 38259 1728
rect 13261 1670 38259 1672
rect 13261 1667 13327 1670
rect 38193 1667 38259 1670
rect 0 1458 800 1488
rect 1393 1458 1459 1461
rect 0 1456 1459 1458
rect 0 1400 1398 1456
rect 1454 1400 1459 1456
rect 0 1398 1459 1400
rect 0 1368 800 1398
rect 1393 1395 1459 1398
rect 2630 1260 2636 1324
rect 2700 1322 2706 1324
rect 34697 1322 34763 1325
rect 2700 1320 34763 1322
rect 2700 1264 34702 1320
rect 34758 1264 34763 1320
rect 2700 1262 34763 1264
rect 2700 1260 2706 1262
rect 34697 1259 34763 1262
rect 39389 98 39455 101
rect 39566 98 40366 128
rect 39389 96 40366 98
rect 39389 40 39394 96
rect 39450 40 40366 96
rect 39389 38 40366 40
rect 39389 35 39455 38
rect 39566 8 40366 38
<< via3 >>
rect 5713 26684 5777 26688
rect 5713 26628 5717 26684
rect 5717 26628 5773 26684
rect 5773 26628 5777 26684
rect 5713 26624 5777 26628
rect 5793 26684 5857 26688
rect 5793 26628 5797 26684
rect 5797 26628 5853 26684
rect 5853 26628 5857 26684
rect 5793 26624 5857 26628
rect 5873 26684 5937 26688
rect 5873 26628 5877 26684
rect 5877 26628 5933 26684
rect 5933 26628 5937 26684
rect 5873 26624 5937 26628
rect 5953 26684 6017 26688
rect 5953 26628 5957 26684
rect 5957 26628 6013 26684
rect 6013 26628 6017 26684
rect 5953 26624 6017 26628
rect 15235 26684 15299 26688
rect 15235 26628 15239 26684
rect 15239 26628 15295 26684
rect 15295 26628 15299 26684
rect 15235 26624 15299 26628
rect 15315 26684 15379 26688
rect 15315 26628 15319 26684
rect 15319 26628 15375 26684
rect 15375 26628 15379 26684
rect 15315 26624 15379 26628
rect 15395 26684 15459 26688
rect 15395 26628 15399 26684
rect 15399 26628 15455 26684
rect 15455 26628 15459 26684
rect 15395 26624 15459 26628
rect 15475 26684 15539 26688
rect 15475 26628 15479 26684
rect 15479 26628 15535 26684
rect 15535 26628 15539 26684
rect 15475 26624 15539 26628
rect 24757 26684 24821 26688
rect 24757 26628 24761 26684
rect 24761 26628 24817 26684
rect 24817 26628 24821 26684
rect 24757 26624 24821 26628
rect 24837 26684 24901 26688
rect 24837 26628 24841 26684
rect 24841 26628 24897 26684
rect 24897 26628 24901 26684
rect 24837 26624 24901 26628
rect 24917 26684 24981 26688
rect 24917 26628 24921 26684
rect 24921 26628 24977 26684
rect 24977 26628 24981 26684
rect 24917 26624 24981 26628
rect 24997 26684 25061 26688
rect 24997 26628 25001 26684
rect 25001 26628 25057 26684
rect 25057 26628 25061 26684
rect 24997 26624 25061 26628
rect 34279 26684 34343 26688
rect 34279 26628 34283 26684
rect 34283 26628 34339 26684
rect 34339 26628 34343 26684
rect 34279 26624 34343 26628
rect 34359 26684 34423 26688
rect 34359 26628 34363 26684
rect 34363 26628 34419 26684
rect 34419 26628 34423 26684
rect 34359 26624 34423 26628
rect 34439 26684 34503 26688
rect 34439 26628 34443 26684
rect 34443 26628 34499 26684
rect 34499 26628 34503 26684
rect 34439 26624 34503 26628
rect 34519 26684 34583 26688
rect 34519 26628 34523 26684
rect 34523 26628 34579 26684
rect 34579 26628 34583 26684
rect 34519 26624 34583 26628
rect 12020 26420 12084 26484
rect 6316 26284 6380 26348
rect 14780 26284 14844 26348
rect 18644 26284 18708 26348
rect 10474 26140 10538 26144
rect 10474 26084 10478 26140
rect 10478 26084 10534 26140
rect 10534 26084 10538 26140
rect 10474 26080 10538 26084
rect 10554 26140 10618 26144
rect 10554 26084 10558 26140
rect 10558 26084 10614 26140
rect 10614 26084 10618 26140
rect 10554 26080 10618 26084
rect 10634 26140 10698 26144
rect 10634 26084 10638 26140
rect 10638 26084 10694 26140
rect 10694 26084 10698 26140
rect 10634 26080 10698 26084
rect 10714 26140 10778 26144
rect 10714 26084 10718 26140
rect 10718 26084 10774 26140
rect 10774 26084 10778 26140
rect 10714 26080 10778 26084
rect 19996 26140 20060 26144
rect 19996 26084 20000 26140
rect 20000 26084 20056 26140
rect 20056 26084 20060 26140
rect 19996 26080 20060 26084
rect 20076 26140 20140 26144
rect 20076 26084 20080 26140
rect 20080 26084 20136 26140
rect 20136 26084 20140 26140
rect 20076 26080 20140 26084
rect 20156 26140 20220 26144
rect 20156 26084 20160 26140
rect 20160 26084 20216 26140
rect 20216 26084 20220 26140
rect 20156 26080 20220 26084
rect 20236 26140 20300 26144
rect 20236 26084 20240 26140
rect 20240 26084 20296 26140
rect 20296 26084 20300 26140
rect 20236 26080 20300 26084
rect 29518 26140 29582 26144
rect 29518 26084 29522 26140
rect 29522 26084 29578 26140
rect 29578 26084 29582 26140
rect 29518 26080 29582 26084
rect 29598 26140 29662 26144
rect 29598 26084 29602 26140
rect 29602 26084 29658 26140
rect 29658 26084 29662 26140
rect 29598 26080 29662 26084
rect 29678 26140 29742 26144
rect 29678 26084 29682 26140
rect 29682 26084 29738 26140
rect 29738 26084 29742 26140
rect 29678 26080 29742 26084
rect 29758 26140 29822 26144
rect 29758 26084 29762 26140
rect 29762 26084 29818 26140
rect 29818 26084 29822 26140
rect 29758 26080 29822 26084
rect 39040 26140 39104 26144
rect 39040 26084 39044 26140
rect 39044 26084 39100 26140
rect 39100 26084 39104 26140
rect 39040 26080 39104 26084
rect 39120 26140 39184 26144
rect 39120 26084 39124 26140
rect 39124 26084 39180 26140
rect 39180 26084 39184 26140
rect 39120 26080 39184 26084
rect 39200 26140 39264 26144
rect 39200 26084 39204 26140
rect 39204 26084 39260 26140
rect 39260 26084 39264 26140
rect 39200 26080 39264 26084
rect 39280 26140 39344 26144
rect 39280 26084 39284 26140
rect 39284 26084 39340 26140
rect 39340 26084 39344 26140
rect 39280 26080 39344 26084
rect 5713 25596 5777 25600
rect 5713 25540 5717 25596
rect 5717 25540 5773 25596
rect 5773 25540 5777 25596
rect 5713 25536 5777 25540
rect 5793 25596 5857 25600
rect 5793 25540 5797 25596
rect 5797 25540 5853 25596
rect 5853 25540 5857 25596
rect 5793 25536 5857 25540
rect 5873 25596 5937 25600
rect 5873 25540 5877 25596
rect 5877 25540 5933 25596
rect 5933 25540 5937 25596
rect 5873 25536 5937 25540
rect 5953 25596 6017 25600
rect 5953 25540 5957 25596
rect 5957 25540 6013 25596
rect 6013 25540 6017 25596
rect 5953 25536 6017 25540
rect 15235 25596 15299 25600
rect 15235 25540 15239 25596
rect 15239 25540 15295 25596
rect 15295 25540 15299 25596
rect 15235 25536 15299 25540
rect 15315 25596 15379 25600
rect 15315 25540 15319 25596
rect 15319 25540 15375 25596
rect 15375 25540 15379 25596
rect 15315 25536 15379 25540
rect 15395 25596 15459 25600
rect 15395 25540 15399 25596
rect 15399 25540 15455 25596
rect 15455 25540 15459 25596
rect 15395 25536 15459 25540
rect 15475 25596 15539 25600
rect 15475 25540 15479 25596
rect 15479 25540 15535 25596
rect 15535 25540 15539 25596
rect 15475 25536 15539 25540
rect 24757 25596 24821 25600
rect 24757 25540 24761 25596
rect 24761 25540 24817 25596
rect 24817 25540 24821 25596
rect 24757 25536 24821 25540
rect 24837 25596 24901 25600
rect 24837 25540 24841 25596
rect 24841 25540 24897 25596
rect 24897 25540 24901 25596
rect 24837 25536 24901 25540
rect 24917 25596 24981 25600
rect 24917 25540 24921 25596
rect 24921 25540 24977 25596
rect 24977 25540 24981 25596
rect 24917 25536 24981 25540
rect 24997 25596 25061 25600
rect 24997 25540 25001 25596
rect 25001 25540 25057 25596
rect 25057 25540 25061 25596
rect 24997 25536 25061 25540
rect 34279 25596 34343 25600
rect 34279 25540 34283 25596
rect 34283 25540 34339 25596
rect 34339 25540 34343 25596
rect 34279 25536 34343 25540
rect 34359 25596 34423 25600
rect 34359 25540 34363 25596
rect 34363 25540 34419 25596
rect 34419 25540 34423 25596
rect 34359 25536 34423 25540
rect 34439 25596 34503 25600
rect 34439 25540 34443 25596
rect 34443 25540 34499 25596
rect 34499 25540 34503 25596
rect 34439 25536 34503 25540
rect 34519 25596 34583 25600
rect 34519 25540 34523 25596
rect 34523 25540 34579 25596
rect 34579 25540 34583 25596
rect 34519 25536 34583 25540
rect 23980 25196 24044 25260
rect 10474 25052 10538 25056
rect 10474 24996 10478 25052
rect 10478 24996 10534 25052
rect 10534 24996 10538 25052
rect 10474 24992 10538 24996
rect 10554 25052 10618 25056
rect 10554 24996 10558 25052
rect 10558 24996 10614 25052
rect 10614 24996 10618 25052
rect 10554 24992 10618 24996
rect 10634 25052 10698 25056
rect 10634 24996 10638 25052
rect 10638 24996 10694 25052
rect 10694 24996 10698 25052
rect 10634 24992 10698 24996
rect 10714 25052 10778 25056
rect 10714 24996 10718 25052
rect 10718 24996 10774 25052
rect 10774 24996 10778 25052
rect 10714 24992 10778 24996
rect 19996 25052 20060 25056
rect 19996 24996 20000 25052
rect 20000 24996 20056 25052
rect 20056 24996 20060 25052
rect 19996 24992 20060 24996
rect 20076 25052 20140 25056
rect 20076 24996 20080 25052
rect 20080 24996 20136 25052
rect 20136 24996 20140 25052
rect 20076 24992 20140 24996
rect 20156 25052 20220 25056
rect 20156 24996 20160 25052
rect 20160 24996 20216 25052
rect 20216 24996 20220 25052
rect 20156 24992 20220 24996
rect 20236 25052 20300 25056
rect 20236 24996 20240 25052
rect 20240 24996 20296 25052
rect 20296 24996 20300 25052
rect 20236 24992 20300 24996
rect 29518 25052 29582 25056
rect 29518 24996 29522 25052
rect 29522 24996 29578 25052
rect 29578 24996 29582 25052
rect 29518 24992 29582 24996
rect 29598 25052 29662 25056
rect 29598 24996 29602 25052
rect 29602 24996 29658 25052
rect 29658 24996 29662 25052
rect 29598 24992 29662 24996
rect 29678 25052 29742 25056
rect 29678 24996 29682 25052
rect 29682 24996 29738 25052
rect 29738 24996 29742 25052
rect 29678 24992 29742 24996
rect 29758 25052 29822 25056
rect 29758 24996 29762 25052
rect 29762 24996 29818 25052
rect 29818 24996 29822 25052
rect 29758 24992 29822 24996
rect 39040 25052 39104 25056
rect 39040 24996 39044 25052
rect 39044 24996 39100 25052
rect 39100 24996 39104 25052
rect 39040 24992 39104 24996
rect 39120 25052 39184 25056
rect 39120 24996 39124 25052
rect 39124 24996 39180 25052
rect 39180 24996 39184 25052
rect 39120 24992 39184 24996
rect 39200 25052 39264 25056
rect 39200 24996 39204 25052
rect 39204 24996 39260 25052
rect 39260 24996 39264 25052
rect 39200 24992 39264 24996
rect 39280 25052 39344 25056
rect 39280 24996 39284 25052
rect 39284 24996 39340 25052
rect 39340 24996 39344 25052
rect 39280 24992 39344 24996
rect 13124 24712 13188 24716
rect 13124 24656 13138 24712
rect 13138 24656 13188 24712
rect 13124 24652 13188 24656
rect 16620 24652 16684 24716
rect 5713 24508 5777 24512
rect 5713 24452 5717 24508
rect 5717 24452 5773 24508
rect 5773 24452 5777 24508
rect 5713 24448 5777 24452
rect 5793 24508 5857 24512
rect 5793 24452 5797 24508
rect 5797 24452 5853 24508
rect 5853 24452 5857 24508
rect 5793 24448 5857 24452
rect 5873 24508 5937 24512
rect 5873 24452 5877 24508
rect 5877 24452 5933 24508
rect 5933 24452 5937 24508
rect 5873 24448 5937 24452
rect 5953 24508 6017 24512
rect 5953 24452 5957 24508
rect 5957 24452 6013 24508
rect 6013 24452 6017 24508
rect 5953 24448 6017 24452
rect 15235 24508 15299 24512
rect 15235 24452 15239 24508
rect 15239 24452 15295 24508
rect 15295 24452 15299 24508
rect 15235 24448 15299 24452
rect 15315 24508 15379 24512
rect 15315 24452 15319 24508
rect 15319 24452 15375 24508
rect 15375 24452 15379 24508
rect 15315 24448 15379 24452
rect 15395 24508 15459 24512
rect 15395 24452 15399 24508
rect 15399 24452 15455 24508
rect 15455 24452 15459 24508
rect 15395 24448 15459 24452
rect 15475 24508 15539 24512
rect 15475 24452 15479 24508
rect 15479 24452 15535 24508
rect 15535 24452 15539 24508
rect 15475 24448 15539 24452
rect 24757 24508 24821 24512
rect 24757 24452 24761 24508
rect 24761 24452 24817 24508
rect 24817 24452 24821 24508
rect 24757 24448 24821 24452
rect 24837 24508 24901 24512
rect 24837 24452 24841 24508
rect 24841 24452 24897 24508
rect 24897 24452 24901 24508
rect 24837 24448 24901 24452
rect 24917 24508 24981 24512
rect 24917 24452 24921 24508
rect 24921 24452 24977 24508
rect 24977 24452 24981 24508
rect 24917 24448 24981 24452
rect 24997 24508 25061 24512
rect 24997 24452 25001 24508
rect 25001 24452 25057 24508
rect 25057 24452 25061 24508
rect 24997 24448 25061 24452
rect 34279 24508 34343 24512
rect 34279 24452 34283 24508
rect 34283 24452 34339 24508
rect 34339 24452 34343 24508
rect 34279 24448 34343 24452
rect 34359 24508 34423 24512
rect 34359 24452 34363 24508
rect 34363 24452 34419 24508
rect 34419 24452 34423 24508
rect 34359 24448 34423 24452
rect 34439 24508 34503 24512
rect 34439 24452 34443 24508
rect 34443 24452 34499 24508
rect 34499 24452 34503 24508
rect 34439 24448 34503 24452
rect 34519 24508 34583 24512
rect 34519 24452 34523 24508
rect 34523 24452 34579 24508
rect 34579 24452 34583 24508
rect 34519 24448 34583 24452
rect 17172 24108 17236 24172
rect 10474 23964 10538 23968
rect 10474 23908 10478 23964
rect 10478 23908 10534 23964
rect 10534 23908 10538 23964
rect 10474 23904 10538 23908
rect 10554 23964 10618 23968
rect 10554 23908 10558 23964
rect 10558 23908 10614 23964
rect 10614 23908 10618 23964
rect 10554 23904 10618 23908
rect 10634 23964 10698 23968
rect 10634 23908 10638 23964
rect 10638 23908 10694 23964
rect 10694 23908 10698 23964
rect 10634 23904 10698 23908
rect 10714 23964 10778 23968
rect 10714 23908 10718 23964
rect 10718 23908 10774 23964
rect 10774 23908 10778 23964
rect 10714 23904 10778 23908
rect 19996 23964 20060 23968
rect 19996 23908 20000 23964
rect 20000 23908 20056 23964
rect 20056 23908 20060 23964
rect 19996 23904 20060 23908
rect 20076 23964 20140 23968
rect 20076 23908 20080 23964
rect 20080 23908 20136 23964
rect 20136 23908 20140 23964
rect 20076 23904 20140 23908
rect 20156 23964 20220 23968
rect 20156 23908 20160 23964
rect 20160 23908 20216 23964
rect 20216 23908 20220 23964
rect 20156 23904 20220 23908
rect 20236 23964 20300 23968
rect 20236 23908 20240 23964
rect 20240 23908 20296 23964
rect 20296 23908 20300 23964
rect 20236 23904 20300 23908
rect 29518 23964 29582 23968
rect 29518 23908 29522 23964
rect 29522 23908 29578 23964
rect 29578 23908 29582 23964
rect 29518 23904 29582 23908
rect 29598 23964 29662 23968
rect 29598 23908 29602 23964
rect 29602 23908 29658 23964
rect 29658 23908 29662 23964
rect 29598 23904 29662 23908
rect 29678 23964 29742 23968
rect 29678 23908 29682 23964
rect 29682 23908 29738 23964
rect 29738 23908 29742 23964
rect 29678 23904 29742 23908
rect 29758 23964 29822 23968
rect 29758 23908 29762 23964
rect 29762 23908 29818 23964
rect 29818 23908 29822 23964
rect 29758 23904 29822 23908
rect 39040 23964 39104 23968
rect 39040 23908 39044 23964
rect 39044 23908 39100 23964
rect 39100 23908 39104 23964
rect 39040 23904 39104 23908
rect 39120 23964 39184 23968
rect 39120 23908 39124 23964
rect 39124 23908 39180 23964
rect 39180 23908 39184 23964
rect 39120 23904 39184 23908
rect 39200 23964 39264 23968
rect 39200 23908 39204 23964
rect 39204 23908 39260 23964
rect 39260 23908 39264 23964
rect 39200 23904 39264 23908
rect 39280 23964 39344 23968
rect 39280 23908 39284 23964
rect 39284 23908 39340 23964
rect 39340 23908 39344 23964
rect 39280 23904 39344 23908
rect 18828 23428 18892 23492
rect 5713 23420 5777 23424
rect 5713 23364 5717 23420
rect 5717 23364 5773 23420
rect 5773 23364 5777 23420
rect 5713 23360 5777 23364
rect 5793 23420 5857 23424
rect 5793 23364 5797 23420
rect 5797 23364 5853 23420
rect 5853 23364 5857 23420
rect 5793 23360 5857 23364
rect 5873 23420 5937 23424
rect 5873 23364 5877 23420
rect 5877 23364 5933 23420
rect 5933 23364 5937 23420
rect 5873 23360 5937 23364
rect 5953 23420 6017 23424
rect 5953 23364 5957 23420
rect 5957 23364 6013 23420
rect 6013 23364 6017 23420
rect 5953 23360 6017 23364
rect 15235 23420 15299 23424
rect 15235 23364 15239 23420
rect 15239 23364 15295 23420
rect 15295 23364 15299 23420
rect 15235 23360 15299 23364
rect 15315 23420 15379 23424
rect 15315 23364 15319 23420
rect 15319 23364 15375 23420
rect 15375 23364 15379 23420
rect 15315 23360 15379 23364
rect 15395 23420 15459 23424
rect 15395 23364 15399 23420
rect 15399 23364 15455 23420
rect 15455 23364 15459 23420
rect 15395 23360 15459 23364
rect 15475 23420 15539 23424
rect 15475 23364 15479 23420
rect 15479 23364 15535 23420
rect 15535 23364 15539 23420
rect 15475 23360 15539 23364
rect 24757 23420 24821 23424
rect 24757 23364 24761 23420
rect 24761 23364 24817 23420
rect 24817 23364 24821 23420
rect 24757 23360 24821 23364
rect 24837 23420 24901 23424
rect 24837 23364 24841 23420
rect 24841 23364 24897 23420
rect 24897 23364 24901 23420
rect 24837 23360 24901 23364
rect 24917 23420 24981 23424
rect 24917 23364 24921 23420
rect 24921 23364 24977 23420
rect 24977 23364 24981 23420
rect 24917 23360 24981 23364
rect 24997 23420 25061 23424
rect 24997 23364 25001 23420
rect 25001 23364 25057 23420
rect 25057 23364 25061 23420
rect 24997 23360 25061 23364
rect 34279 23420 34343 23424
rect 34279 23364 34283 23420
rect 34283 23364 34339 23420
rect 34339 23364 34343 23420
rect 34279 23360 34343 23364
rect 34359 23420 34423 23424
rect 34359 23364 34363 23420
rect 34363 23364 34419 23420
rect 34419 23364 34423 23420
rect 34359 23360 34423 23364
rect 34439 23420 34503 23424
rect 34439 23364 34443 23420
rect 34443 23364 34499 23420
rect 34499 23364 34503 23420
rect 34439 23360 34503 23364
rect 34519 23420 34583 23424
rect 34519 23364 34523 23420
rect 34523 23364 34579 23420
rect 34579 23364 34583 23420
rect 34519 23360 34583 23364
rect 25636 22884 25700 22948
rect 10474 22876 10538 22880
rect 10474 22820 10478 22876
rect 10478 22820 10534 22876
rect 10534 22820 10538 22876
rect 10474 22816 10538 22820
rect 10554 22876 10618 22880
rect 10554 22820 10558 22876
rect 10558 22820 10614 22876
rect 10614 22820 10618 22876
rect 10554 22816 10618 22820
rect 10634 22876 10698 22880
rect 10634 22820 10638 22876
rect 10638 22820 10694 22876
rect 10694 22820 10698 22876
rect 10634 22816 10698 22820
rect 10714 22876 10778 22880
rect 10714 22820 10718 22876
rect 10718 22820 10774 22876
rect 10774 22820 10778 22876
rect 10714 22816 10778 22820
rect 19996 22876 20060 22880
rect 19996 22820 20000 22876
rect 20000 22820 20056 22876
rect 20056 22820 20060 22876
rect 19996 22816 20060 22820
rect 20076 22876 20140 22880
rect 20076 22820 20080 22876
rect 20080 22820 20136 22876
rect 20136 22820 20140 22876
rect 20076 22816 20140 22820
rect 20156 22876 20220 22880
rect 20156 22820 20160 22876
rect 20160 22820 20216 22876
rect 20216 22820 20220 22876
rect 20156 22816 20220 22820
rect 20236 22876 20300 22880
rect 20236 22820 20240 22876
rect 20240 22820 20296 22876
rect 20296 22820 20300 22876
rect 20236 22816 20300 22820
rect 29518 22876 29582 22880
rect 29518 22820 29522 22876
rect 29522 22820 29578 22876
rect 29578 22820 29582 22876
rect 29518 22816 29582 22820
rect 29598 22876 29662 22880
rect 29598 22820 29602 22876
rect 29602 22820 29658 22876
rect 29658 22820 29662 22876
rect 29598 22816 29662 22820
rect 29678 22876 29742 22880
rect 29678 22820 29682 22876
rect 29682 22820 29738 22876
rect 29738 22820 29742 22876
rect 29678 22816 29742 22820
rect 29758 22876 29822 22880
rect 29758 22820 29762 22876
rect 29762 22820 29818 22876
rect 29818 22820 29822 22876
rect 29758 22816 29822 22820
rect 39040 22876 39104 22880
rect 39040 22820 39044 22876
rect 39044 22820 39100 22876
rect 39100 22820 39104 22876
rect 39040 22816 39104 22820
rect 39120 22876 39184 22880
rect 39120 22820 39124 22876
rect 39124 22820 39180 22876
rect 39180 22820 39184 22876
rect 39120 22816 39184 22820
rect 39200 22876 39264 22880
rect 39200 22820 39204 22876
rect 39204 22820 39260 22876
rect 39260 22820 39264 22876
rect 39200 22816 39264 22820
rect 39280 22876 39344 22880
rect 39280 22820 39284 22876
rect 39284 22820 39340 22876
rect 39340 22820 39344 22876
rect 39280 22816 39344 22820
rect 30236 22340 30300 22404
rect 5713 22332 5777 22336
rect 5713 22276 5717 22332
rect 5717 22276 5773 22332
rect 5773 22276 5777 22332
rect 5713 22272 5777 22276
rect 5793 22332 5857 22336
rect 5793 22276 5797 22332
rect 5797 22276 5853 22332
rect 5853 22276 5857 22332
rect 5793 22272 5857 22276
rect 5873 22332 5937 22336
rect 5873 22276 5877 22332
rect 5877 22276 5933 22332
rect 5933 22276 5937 22332
rect 5873 22272 5937 22276
rect 5953 22332 6017 22336
rect 5953 22276 5957 22332
rect 5957 22276 6013 22332
rect 6013 22276 6017 22332
rect 5953 22272 6017 22276
rect 15235 22332 15299 22336
rect 15235 22276 15239 22332
rect 15239 22276 15295 22332
rect 15295 22276 15299 22332
rect 15235 22272 15299 22276
rect 15315 22332 15379 22336
rect 15315 22276 15319 22332
rect 15319 22276 15375 22332
rect 15375 22276 15379 22332
rect 15315 22272 15379 22276
rect 15395 22332 15459 22336
rect 15395 22276 15399 22332
rect 15399 22276 15455 22332
rect 15455 22276 15459 22332
rect 15395 22272 15459 22276
rect 15475 22332 15539 22336
rect 15475 22276 15479 22332
rect 15479 22276 15535 22332
rect 15535 22276 15539 22332
rect 15475 22272 15539 22276
rect 24757 22332 24821 22336
rect 24757 22276 24761 22332
rect 24761 22276 24817 22332
rect 24817 22276 24821 22332
rect 24757 22272 24821 22276
rect 24837 22332 24901 22336
rect 24837 22276 24841 22332
rect 24841 22276 24897 22332
rect 24897 22276 24901 22332
rect 24837 22272 24901 22276
rect 24917 22332 24981 22336
rect 24917 22276 24921 22332
rect 24921 22276 24977 22332
rect 24977 22276 24981 22332
rect 24917 22272 24981 22276
rect 24997 22332 25061 22336
rect 24997 22276 25001 22332
rect 25001 22276 25057 22332
rect 25057 22276 25061 22332
rect 24997 22272 25061 22276
rect 34279 22332 34343 22336
rect 34279 22276 34283 22332
rect 34283 22276 34339 22332
rect 34339 22276 34343 22332
rect 34279 22272 34343 22276
rect 34359 22332 34423 22336
rect 34359 22276 34363 22332
rect 34363 22276 34419 22332
rect 34419 22276 34423 22332
rect 34359 22272 34423 22276
rect 34439 22332 34503 22336
rect 34439 22276 34443 22332
rect 34443 22276 34499 22332
rect 34499 22276 34503 22332
rect 34439 22272 34503 22276
rect 34519 22332 34583 22336
rect 34519 22276 34523 22332
rect 34523 22276 34579 22332
rect 34579 22276 34583 22332
rect 34519 22272 34583 22276
rect 33180 22068 33244 22132
rect 32996 21796 33060 21860
rect 10474 21788 10538 21792
rect 10474 21732 10478 21788
rect 10478 21732 10534 21788
rect 10534 21732 10538 21788
rect 10474 21728 10538 21732
rect 10554 21788 10618 21792
rect 10554 21732 10558 21788
rect 10558 21732 10614 21788
rect 10614 21732 10618 21788
rect 10554 21728 10618 21732
rect 10634 21788 10698 21792
rect 10634 21732 10638 21788
rect 10638 21732 10694 21788
rect 10694 21732 10698 21788
rect 10634 21728 10698 21732
rect 10714 21788 10778 21792
rect 10714 21732 10718 21788
rect 10718 21732 10774 21788
rect 10774 21732 10778 21788
rect 10714 21728 10778 21732
rect 19996 21788 20060 21792
rect 19996 21732 20000 21788
rect 20000 21732 20056 21788
rect 20056 21732 20060 21788
rect 19996 21728 20060 21732
rect 20076 21788 20140 21792
rect 20076 21732 20080 21788
rect 20080 21732 20136 21788
rect 20136 21732 20140 21788
rect 20076 21728 20140 21732
rect 20156 21788 20220 21792
rect 20156 21732 20160 21788
rect 20160 21732 20216 21788
rect 20216 21732 20220 21788
rect 20156 21728 20220 21732
rect 20236 21788 20300 21792
rect 20236 21732 20240 21788
rect 20240 21732 20296 21788
rect 20296 21732 20300 21788
rect 20236 21728 20300 21732
rect 29518 21788 29582 21792
rect 29518 21732 29522 21788
rect 29522 21732 29578 21788
rect 29578 21732 29582 21788
rect 29518 21728 29582 21732
rect 29598 21788 29662 21792
rect 29598 21732 29602 21788
rect 29602 21732 29658 21788
rect 29658 21732 29662 21788
rect 29598 21728 29662 21732
rect 29678 21788 29742 21792
rect 29678 21732 29682 21788
rect 29682 21732 29738 21788
rect 29738 21732 29742 21788
rect 29678 21728 29742 21732
rect 29758 21788 29822 21792
rect 29758 21732 29762 21788
rect 29762 21732 29818 21788
rect 29818 21732 29822 21788
rect 29758 21728 29822 21732
rect 39040 21788 39104 21792
rect 39040 21732 39044 21788
rect 39044 21732 39100 21788
rect 39100 21732 39104 21788
rect 39040 21728 39104 21732
rect 39120 21788 39184 21792
rect 39120 21732 39124 21788
rect 39124 21732 39180 21788
rect 39180 21732 39184 21788
rect 39120 21728 39184 21732
rect 39200 21788 39264 21792
rect 39200 21732 39204 21788
rect 39204 21732 39260 21788
rect 39260 21732 39264 21788
rect 39200 21728 39264 21732
rect 39280 21788 39344 21792
rect 39280 21732 39284 21788
rect 39284 21732 39340 21788
rect 39340 21732 39344 21788
rect 39280 21728 39344 21732
rect 5713 21244 5777 21248
rect 5713 21188 5717 21244
rect 5717 21188 5773 21244
rect 5773 21188 5777 21244
rect 5713 21184 5777 21188
rect 5793 21244 5857 21248
rect 5793 21188 5797 21244
rect 5797 21188 5853 21244
rect 5853 21188 5857 21244
rect 5793 21184 5857 21188
rect 5873 21244 5937 21248
rect 5873 21188 5877 21244
rect 5877 21188 5933 21244
rect 5933 21188 5937 21244
rect 5873 21184 5937 21188
rect 5953 21244 6017 21248
rect 5953 21188 5957 21244
rect 5957 21188 6013 21244
rect 6013 21188 6017 21244
rect 5953 21184 6017 21188
rect 15235 21244 15299 21248
rect 15235 21188 15239 21244
rect 15239 21188 15295 21244
rect 15295 21188 15299 21244
rect 15235 21184 15299 21188
rect 15315 21244 15379 21248
rect 15315 21188 15319 21244
rect 15319 21188 15375 21244
rect 15375 21188 15379 21244
rect 15315 21184 15379 21188
rect 15395 21244 15459 21248
rect 15395 21188 15399 21244
rect 15399 21188 15455 21244
rect 15455 21188 15459 21244
rect 15395 21184 15459 21188
rect 15475 21244 15539 21248
rect 15475 21188 15479 21244
rect 15479 21188 15535 21244
rect 15535 21188 15539 21244
rect 15475 21184 15539 21188
rect 24757 21244 24821 21248
rect 24757 21188 24761 21244
rect 24761 21188 24817 21244
rect 24817 21188 24821 21244
rect 24757 21184 24821 21188
rect 24837 21244 24901 21248
rect 24837 21188 24841 21244
rect 24841 21188 24897 21244
rect 24897 21188 24901 21244
rect 24837 21184 24901 21188
rect 24917 21244 24981 21248
rect 24917 21188 24921 21244
rect 24921 21188 24977 21244
rect 24977 21188 24981 21244
rect 24917 21184 24981 21188
rect 24997 21244 25061 21248
rect 24997 21188 25001 21244
rect 25001 21188 25057 21244
rect 25057 21188 25061 21244
rect 24997 21184 25061 21188
rect 34279 21244 34343 21248
rect 34279 21188 34283 21244
rect 34283 21188 34339 21244
rect 34339 21188 34343 21244
rect 34279 21184 34343 21188
rect 34359 21244 34423 21248
rect 34359 21188 34363 21244
rect 34363 21188 34419 21244
rect 34419 21188 34423 21244
rect 34359 21184 34423 21188
rect 34439 21244 34503 21248
rect 34439 21188 34443 21244
rect 34443 21188 34499 21244
rect 34499 21188 34503 21244
rect 34439 21184 34503 21188
rect 34519 21244 34583 21248
rect 34519 21188 34523 21244
rect 34523 21188 34579 21244
rect 34579 21188 34583 21244
rect 34519 21184 34583 21188
rect 22692 20980 22756 21044
rect 12756 20844 12820 20908
rect 17908 20708 17972 20772
rect 32812 20768 32876 20772
rect 32812 20712 32826 20768
rect 32826 20712 32876 20768
rect 32812 20708 32876 20712
rect 10474 20700 10538 20704
rect 10474 20644 10478 20700
rect 10478 20644 10534 20700
rect 10534 20644 10538 20700
rect 10474 20640 10538 20644
rect 10554 20700 10618 20704
rect 10554 20644 10558 20700
rect 10558 20644 10614 20700
rect 10614 20644 10618 20700
rect 10554 20640 10618 20644
rect 10634 20700 10698 20704
rect 10634 20644 10638 20700
rect 10638 20644 10694 20700
rect 10694 20644 10698 20700
rect 10634 20640 10698 20644
rect 10714 20700 10778 20704
rect 10714 20644 10718 20700
rect 10718 20644 10774 20700
rect 10774 20644 10778 20700
rect 10714 20640 10778 20644
rect 19996 20700 20060 20704
rect 19996 20644 20000 20700
rect 20000 20644 20056 20700
rect 20056 20644 20060 20700
rect 19996 20640 20060 20644
rect 20076 20700 20140 20704
rect 20076 20644 20080 20700
rect 20080 20644 20136 20700
rect 20136 20644 20140 20700
rect 20076 20640 20140 20644
rect 20156 20700 20220 20704
rect 20156 20644 20160 20700
rect 20160 20644 20216 20700
rect 20216 20644 20220 20700
rect 20156 20640 20220 20644
rect 20236 20700 20300 20704
rect 20236 20644 20240 20700
rect 20240 20644 20296 20700
rect 20296 20644 20300 20700
rect 20236 20640 20300 20644
rect 29518 20700 29582 20704
rect 29518 20644 29522 20700
rect 29522 20644 29578 20700
rect 29578 20644 29582 20700
rect 29518 20640 29582 20644
rect 29598 20700 29662 20704
rect 29598 20644 29602 20700
rect 29602 20644 29658 20700
rect 29658 20644 29662 20700
rect 29598 20640 29662 20644
rect 29678 20700 29742 20704
rect 29678 20644 29682 20700
rect 29682 20644 29738 20700
rect 29738 20644 29742 20700
rect 29678 20640 29742 20644
rect 29758 20700 29822 20704
rect 29758 20644 29762 20700
rect 29762 20644 29818 20700
rect 29818 20644 29822 20700
rect 29758 20640 29822 20644
rect 39040 20700 39104 20704
rect 39040 20644 39044 20700
rect 39044 20644 39100 20700
rect 39100 20644 39104 20700
rect 39040 20640 39104 20644
rect 39120 20700 39184 20704
rect 39120 20644 39124 20700
rect 39124 20644 39180 20700
rect 39180 20644 39184 20700
rect 39120 20640 39184 20644
rect 39200 20700 39264 20704
rect 39200 20644 39204 20700
rect 39204 20644 39260 20700
rect 39260 20644 39264 20700
rect 39200 20640 39264 20644
rect 39280 20700 39344 20704
rect 39280 20644 39284 20700
rect 39284 20644 39340 20700
rect 39340 20644 39344 20700
rect 39280 20640 39344 20644
rect 5713 20156 5777 20160
rect 5713 20100 5717 20156
rect 5717 20100 5773 20156
rect 5773 20100 5777 20156
rect 5713 20096 5777 20100
rect 5793 20156 5857 20160
rect 5793 20100 5797 20156
rect 5797 20100 5853 20156
rect 5853 20100 5857 20156
rect 5793 20096 5857 20100
rect 5873 20156 5937 20160
rect 5873 20100 5877 20156
rect 5877 20100 5933 20156
rect 5933 20100 5937 20156
rect 5873 20096 5937 20100
rect 5953 20156 6017 20160
rect 5953 20100 5957 20156
rect 5957 20100 6013 20156
rect 6013 20100 6017 20156
rect 5953 20096 6017 20100
rect 15235 20156 15299 20160
rect 15235 20100 15239 20156
rect 15239 20100 15295 20156
rect 15295 20100 15299 20156
rect 15235 20096 15299 20100
rect 15315 20156 15379 20160
rect 15315 20100 15319 20156
rect 15319 20100 15375 20156
rect 15375 20100 15379 20156
rect 15315 20096 15379 20100
rect 15395 20156 15459 20160
rect 15395 20100 15399 20156
rect 15399 20100 15455 20156
rect 15455 20100 15459 20156
rect 15395 20096 15459 20100
rect 15475 20156 15539 20160
rect 15475 20100 15479 20156
rect 15479 20100 15535 20156
rect 15535 20100 15539 20156
rect 15475 20096 15539 20100
rect 24757 20156 24821 20160
rect 24757 20100 24761 20156
rect 24761 20100 24817 20156
rect 24817 20100 24821 20156
rect 24757 20096 24821 20100
rect 24837 20156 24901 20160
rect 24837 20100 24841 20156
rect 24841 20100 24897 20156
rect 24897 20100 24901 20156
rect 24837 20096 24901 20100
rect 24917 20156 24981 20160
rect 24917 20100 24921 20156
rect 24921 20100 24977 20156
rect 24977 20100 24981 20156
rect 24917 20096 24981 20100
rect 24997 20156 25061 20160
rect 24997 20100 25001 20156
rect 25001 20100 25057 20156
rect 25057 20100 25061 20156
rect 24997 20096 25061 20100
rect 34279 20156 34343 20160
rect 34279 20100 34283 20156
rect 34283 20100 34339 20156
rect 34339 20100 34343 20156
rect 34279 20096 34343 20100
rect 34359 20156 34423 20160
rect 34359 20100 34363 20156
rect 34363 20100 34419 20156
rect 34419 20100 34423 20156
rect 34359 20096 34423 20100
rect 34439 20156 34503 20160
rect 34439 20100 34443 20156
rect 34443 20100 34499 20156
rect 34499 20100 34503 20156
rect 34439 20096 34503 20100
rect 34519 20156 34583 20160
rect 34519 20100 34523 20156
rect 34523 20100 34579 20156
rect 34579 20100 34583 20156
rect 34519 20096 34583 20100
rect 14964 19620 15028 19684
rect 10474 19612 10538 19616
rect 10474 19556 10478 19612
rect 10478 19556 10534 19612
rect 10534 19556 10538 19612
rect 10474 19552 10538 19556
rect 10554 19612 10618 19616
rect 10554 19556 10558 19612
rect 10558 19556 10614 19612
rect 10614 19556 10618 19612
rect 10554 19552 10618 19556
rect 10634 19612 10698 19616
rect 10634 19556 10638 19612
rect 10638 19556 10694 19612
rect 10694 19556 10698 19612
rect 10634 19552 10698 19556
rect 10714 19612 10778 19616
rect 10714 19556 10718 19612
rect 10718 19556 10774 19612
rect 10774 19556 10778 19612
rect 10714 19552 10778 19556
rect 19996 19612 20060 19616
rect 19996 19556 20000 19612
rect 20000 19556 20056 19612
rect 20056 19556 20060 19612
rect 19996 19552 20060 19556
rect 20076 19612 20140 19616
rect 20076 19556 20080 19612
rect 20080 19556 20136 19612
rect 20136 19556 20140 19612
rect 20076 19552 20140 19556
rect 20156 19612 20220 19616
rect 20156 19556 20160 19612
rect 20160 19556 20216 19612
rect 20216 19556 20220 19612
rect 20156 19552 20220 19556
rect 20236 19612 20300 19616
rect 20236 19556 20240 19612
rect 20240 19556 20296 19612
rect 20296 19556 20300 19612
rect 20236 19552 20300 19556
rect 29518 19612 29582 19616
rect 29518 19556 29522 19612
rect 29522 19556 29578 19612
rect 29578 19556 29582 19612
rect 29518 19552 29582 19556
rect 29598 19612 29662 19616
rect 29598 19556 29602 19612
rect 29602 19556 29658 19612
rect 29658 19556 29662 19612
rect 29598 19552 29662 19556
rect 29678 19612 29742 19616
rect 29678 19556 29682 19612
rect 29682 19556 29738 19612
rect 29738 19556 29742 19612
rect 29678 19552 29742 19556
rect 29758 19612 29822 19616
rect 29758 19556 29762 19612
rect 29762 19556 29818 19612
rect 29818 19556 29822 19612
rect 29758 19552 29822 19556
rect 39040 19612 39104 19616
rect 39040 19556 39044 19612
rect 39044 19556 39100 19612
rect 39100 19556 39104 19612
rect 39040 19552 39104 19556
rect 39120 19612 39184 19616
rect 39120 19556 39124 19612
rect 39124 19556 39180 19612
rect 39180 19556 39184 19612
rect 39120 19552 39184 19556
rect 39200 19612 39264 19616
rect 39200 19556 39204 19612
rect 39204 19556 39260 19612
rect 39260 19556 39264 19612
rect 39200 19552 39264 19556
rect 39280 19612 39344 19616
rect 39280 19556 39284 19612
rect 39284 19556 39340 19612
rect 39340 19556 39344 19612
rect 39280 19552 39344 19556
rect 13308 19212 13372 19276
rect 14412 19212 14476 19276
rect 32628 19348 32692 19412
rect 5713 19068 5777 19072
rect 5713 19012 5717 19068
rect 5717 19012 5773 19068
rect 5773 19012 5777 19068
rect 5713 19008 5777 19012
rect 5793 19068 5857 19072
rect 5793 19012 5797 19068
rect 5797 19012 5853 19068
rect 5853 19012 5857 19068
rect 5793 19008 5857 19012
rect 5873 19068 5937 19072
rect 5873 19012 5877 19068
rect 5877 19012 5933 19068
rect 5933 19012 5937 19068
rect 5873 19008 5937 19012
rect 5953 19068 6017 19072
rect 5953 19012 5957 19068
rect 5957 19012 6013 19068
rect 6013 19012 6017 19068
rect 5953 19008 6017 19012
rect 15235 19068 15299 19072
rect 15235 19012 15239 19068
rect 15239 19012 15295 19068
rect 15295 19012 15299 19068
rect 15235 19008 15299 19012
rect 15315 19068 15379 19072
rect 15315 19012 15319 19068
rect 15319 19012 15375 19068
rect 15375 19012 15379 19068
rect 15315 19008 15379 19012
rect 15395 19068 15459 19072
rect 15395 19012 15399 19068
rect 15399 19012 15455 19068
rect 15455 19012 15459 19068
rect 15395 19008 15459 19012
rect 15475 19068 15539 19072
rect 15475 19012 15479 19068
rect 15479 19012 15535 19068
rect 15535 19012 15539 19068
rect 15475 19008 15539 19012
rect 24757 19068 24821 19072
rect 24757 19012 24761 19068
rect 24761 19012 24817 19068
rect 24817 19012 24821 19068
rect 24757 19008 24821 19012
rect 24837 19068 24901 19072
rect 24837 19012 24841 19068
rect 24841 19012 24897 19068
rect 24897 19012 24901 19068
rect 24837 19008 24901 19012
rect 24917 19068 24981 19072
rect 24917 19012 24921 19068
rect 24921 19012 24977 19068
rect 24977 19012 24981 19068
rect 24917 19008 24981 19012
rect 24997 19068 25061 19072
rect 24997 19012 25001 19068
rect 25001 19012 25057 19068
rect 25057 19012 25061 19068
rect 24997 19008 25061 19012
rect 34279 19068 34343 19072
rect 34279 19012 34283 19068
rect 34283 19012 34339 19068
rect 34339 19012 34343 19068
rect 34279 19008 34343 19012
rect 34359 19068 34423 19072
rect 34359 19012 34363 19068
rect 34363 19012 34419 19068
rect 34419 19012 34423 19068
rect 34359 19008 34423 19012
rect 34439 19068 34503 19072
rect 34439 19012 34443 19068
rect 34443 19012 34499 19068
rect 34499 19012 34503 19068
rect 34439 19008 34503 19012
rect 34519 19068 34583 19072
rect 34519 19012 34523 19068
rect 34523 19012 34579 19068
rect 34579 19012 34583 19068
rect 34519 19008 34583 19012
rect 15884 18804 15948 18868
rect 16068 18668 16132 18732
rect 25452 18592 25516 18596
rect 25452 18536 25466 18592
rect 25466 18536 25516 18592
rect 25452 18532 25516 18536
rect 10474 18524 10538 18528
rect 10474 18468 10478 18524
rect 10478 18468 10534 18524
rect 10534 18468 10538 18524
rect 10474 18464 10538 18468
rect 10554 18524 10618 18528
rect 10554 18468 10558 18524
rect 10558 18468 10614 18524
rect 10614 18468 10618 18524
rect 10554 18464 10618 18468
rect 10634 18524 10698 18528
rect 10634 18468 10638 18524
rect 10638 18468 10694 18524
rect 10694 18468 10698 18524
rect 10634 18464 10698 18468
rect 10714 18524 10778 18528
rect 10714 18468 10718 18524
rect 10718 18468 10774 18524
rect 10774 18468 10778 18524
rect 10714 18464 10778 18468
rect 19996 18524 20060 18528
rect 19996 18468 20000 18524
rect 20000 18468 20056 18524
rect 20056 18468 20060 18524
rect 19996 18464 20060 18468
rect 20076 18524 20140 18528
rect 20076 18468 20080 18524
rect 20080 18468 20136 18524
rect 20136 18468 20140 18524
rect 20076 18464 20140 18468
rect 20156 18524 20220 18528
rect 20156 18468 20160 18524
rect 20160 18468 20216 18524
rect 20216 18468 20220 18524
rect 20156 18464 20220 18468
rect 20236 18524 20300 18528
rect 20236 18468 20240 18524
rect 20240 18468 20296 18524
rect 20296 18468 20300 18524
rect 20236 18464 20300 18468
rect 29518 18524 29582 18528
rect 29518 18468 29522 18524
rect 29522 18468 29578 18524
rect 29578 18468 29582 18524
rect 29518 18464 29582 18468
rect 29598 18524 29662 18528
rect 29598 18468 29602 18524
rect 29602 18468 29658 18524
rect 29658 18468 29662 18524
rect 29598 18464 29662 18468
rect 29678 18524 29742 18528
rect 29678 18468 29682 18524
rect 29682 18468 29738 18524
rect 29738 18468 29742 18524
rect 29678 18464 29742 18468
rect 29758 18524 29822 18528
rect 29758 18468 29762 18524
rect 29762 18468 29818 18524
rect 29818 18468 29822 18524
rect 29758 18464 29822 18468
rect 39040 18524 39104 18528
rect 39040 18468 39044 18524
rect 39044 18468 39100 18524
rect 39100 18468 39104 18524
rect 39040 18464 39104 18468
rect 39120 18524 39184 18528
rect 39120 18468 39124 18524
rect 39124 18468 39180 18524
rect 39180 18468 39184 18524
rect 39120 18464 39184 18468
rect 39200 18524 39264 18528
rect 39200 18468 39204 18524
rect 39204 18468 39260 18524
rect 39260 18468 39264 18524
rect 39200 18464 39264 18468
rect 39280 18524 39344 18528
rect 39280 18468 39284 18524
rect 39284 18468 39340 18524
rect 39340 18468 39344 18524
rect 39280 18464 39344 18468
rect 22324 18260 22388 18324
rect 16988 18124 17052 18188
rect 17724 18124 17788 18188
rect 33732 18124 33796 18188
rect 27660 17988 27724 18052
rect 5713 17980 5777 17984
rect 5713 17924 5717 17980
rect 5717 17924 5773 17980
rect 5773 17924 5777 17980
rect 5713 17920 5777 17924
rect 5793 17980 5857 17984
rect 5793 17924 5797 17980
rect 5797 17924 5853 17980
rect 5853 17924 5857 17980
rect 5793 17920 5857 17924
rect 5873 17980 5937 17984
rect 5873 17924 5877 17980
rect 5877 17924 5933 17980
rect 5933 17924 5937 17980
rect 5873 17920 5937 17924
rect 5953 17980 6017 17984
rect 5953 17924 5957 17980
rect 5957 17924 6013 17980
rect 6013 17924 6017 17980
rect 5953 17920 6017 17924
rect 15235 17980 15299 17984
rect 15235 17924 15239 17980
rect 15239 17924 15295 17980
rect 15295 17924 15299 17980
rect 15235 17920 15299 17924
rect 15315 17980 15379 17984
rect 15315 17924 15319 17980
rect 15319 17924 15375 17980
rect 15375 17924 15379 17980
rect 15315 17920 15379 17924
rect 15395 17980 15459 17984
rect 15395 17924 15399 17980
rect 15399 17924 15455 17980
rect 15455 17924 15459 17980
rect 15395 17920 15459 17924
rect 15475 17980 15539 17984
rect 15475 17924 15479 17980
rect 15479 17924 15535 17980
rect 15535 17924 15539 17980
rect 15475 17920 15539 17924
rect 24757 17980 24821 17984
rect 24757 17924 24761 17980
rect 24761 17924 24817 17980
rect 24817 17924 24821 17980
rect 24757 17920 24821 17924
rect 24837 17980 24901 17984
rect 24837 17924 24841 17980
rect 24841 17924 24897 17980
rect 24897 17924 24901 17980
rect 24837 17920 24901 17924
rect 24917 17980 24981 17984
rect 24917 17924 24921 17980
rect 24921 17924 24977 17980
rect 24977 17924 24981 17980
rect 24917 17920 24981 17924
rect 24997 17980 25061 17984
rect 24997 17924 25001 17980
rect 25001 17924 25057 17980
rect 25057 17924 25061 17980
rect 24997 17920 25061 17924
rect 34279 17980 34343 17984
rect 34279 17924 34283 17980
rect 34283 17924 34339 17980
rect 34339 17924 34343 17980
rect 34279 17920 34343 17924
rect 34359 17980 34423 17984
rect 34359 17924 34363 17980
rect 34363 17924 34419 17980
rect 34419 17924 34423 17980
rect 34359 17920 34423 17924
rect 34439 17980 34503 17984
rect 34439 17924 34443 17980
rect 34443 17924 34499 17980
rect 34499 17924 34503 17980
rect 34439 17920 34503 17924
rect 34519 17980 34583 17984
rect 34519 17924 34523 17980
rect 34523 17924 34579 17980
rect 34579 17924 34583 17980
rect 34519 17920 34583 17924
rect 27108 17852 27172 17916
rect 18276 17716 18340 17780
rect 10474 17436 10538 17440
rect 10474 17380 10478 17436
rect 10478 17380 10534 17436
rect 10534 17380 10538 17436
rect 10474 17376 10538 17380
rect 10554 17436 10618 17440
rect 10554 17380 10558 17436
rect 10558 17380 10614 17436
rect 10614 17380 10618 17436
rect 10554 17376 10618 17380
rect 10634 17436 10698 17440
rect 10634 17380 10638 17436
rect 10638 17380 10694 17436
rect 10694 17380 10698 17436
rect 10634 17376 10698 17380
rect 10714 17436 10778 17440
rect 10714 17380 10718 17436
rect 10718 17380 10774 17436
rect 10774 17380 10778 17436
rect 10714 17376 10778 17380
rect 19996 17436 20060 17440
rect 19996 17380 20000 17436
rect 20000 17380 20056 17436
rect 20056 17380 20060 17436
rect 19996 17376 20060 17380
rect 20076 17436 20140 17440
rect 20076 17380 20080 17436
rect 20080 17380 20136 17436
rect 20136 17380 20140 17436
rect 20076 17376 20140 17380
rect 20156 17436 20220 17440
rect 20156 17380 20160 17436
rect 20160 17380 20216 17436
rect 20216 17380 20220 17436
rect 20156 17376 20220 17380
rect 20236 17436 20300 17440
rect 20236 17380 20240 17436
rect 20240 17380 20296 17436
rect 20296 17380 20300 17436
rect 20236 17376 20300 17380
rect 29518 17436 29582 17440
rect 29518 17380 29522 17436
rect 29522 17380 29578 17436
rect 29578 17380 29582 17436
rect 29518 17376 29582 17380
rect 29598 17436 29662 17440
rect 29598 17380 29602 17436
rect 29602 17380 29658 17436
rect 29658 17380 29662 17436
rect 29598 17376 29662 17380
rect 29678 17436 29742 17440
rect 29678 17380 29682 17436
rect 29682 17380 29738 17436
rect 29738 17380 29742 17436
rect 29678 17376 29742 17380
rect 29758 17436 29822 17440
rect 29758 17380 29762 17436
rect 29762 17380 29818 17436
rect 29818 17380 29822 17436
rect 29758 17376 29822 17380
rect 39040 17436 39104 17440
rect 39040 17380 39044 17436
rect 39044 17380 39100 17436
rect 39100 17380 39104 17436
rect 39040 17376 39104 17380
rect 39120 17436 39184 17440
rect 39120 17380 39124 17436
rect 39124 17380 39180 17436
rect 39180 17380 39184 17436
rect 39120 17376 39184 17380
rect 39200 17436 39264 17440
rect 39200 17380 39204 17436
rect 39204 17380 39260 17436
rect 39260 17380 39264 17436
rect 39200 17376 39264 17380
rect 39280 17436 39344 17440
rect 39280 17380 39284 17436
rect 39284 17380 39340 17436
rect 39340 17380 39344 17436
rect 39280 17376 39344 17380
rect 19564 17308 19628 17372
rect 6500 17172 6564 17236
rect 5212 17096 5276 17100
rect 5212 17040 5226 17096
rect 5226 17040 5276 17096
rect 5212 17036 5276 17040
rect 31340 17036 31404 17100
rect 5713 16892 5777 16896
rect 5713 16836 5717 16892
rect 5717 16836 5773 16892
rect 5773 16836 5777 16892
rect 5713 16832 5777 16836
rect 5793 16892 5857 16896
rect 5793 16836 5797 16892
rect 5797 16836 5853 16892
rect 5853 16836 5857 16892
rect 5793 16832 5857 16836
rect 5873 16892 5937 16896
rect 5873 16836 5877 16892
rect 5877 16836 5933 16892
rect 5933 16836 5937 16892
rect 5873 16832 5937 16836
rect 5953 16892 6017 16896
rect 5953 16836 5957 16892
rect 5957 16836 6013 16892
rect 6013 16836 6017 16892
rect 5953 16832 6017 16836
rect 15235 16892 15299 16896
rect 15235 16836 15239 16892
rect 15239 16836 15295 16892
rect 15295 16836 15299 16892
rect 15235 16832 15299 16836
rect 15315 16892 15379 16896
rect 15315 16836 15319 16892
rect 15319 16836 15375 16892
rect 15375 16836 15379 16892
rect 15315 16832 15379 16836
rect 15395 16892 15459 16896
rect 15395 16836 15399 16892
rect 15399 16836 15455 16892
rect 15455 16836 15459 16892
rect 15395 16832 15459 16836
rect 15475 16892 15539 16896
rect 15475 16836 15479 16892
rect 15479 16836 15535 16892
rect 15535 16836 15539 16892
rect 15475 16832 15539 16836
rect 24757 16892 24821 16896
rect 24757 16836 24761 16892
rect 24761 16836 24817 16892
rect 24817 16836 24821 16892
rect 24757 16832 24821 16836
rect 24837 16892 24901 16896
rect 24837 16836 24841 16892
rect 24841 16836 24897 16892
rect 24897 16836 24901 16892
rect 24837 16832 24901 16836
rect 24917 16892 24981 16896
rect 24917 16836 24921 16892
rect 24921 16836 24977 16892
rect 24977 16836 24981 16892
rect 24917 16832 24981 16836
rect 24997 16892 25061 16896
rect 24997 16836 25001 16892
rect 25001 16836 25057 16892
rect 25057 16836 25061 16892
rect 24997 16832 25061 16836
rect 34279 16892 34343 16896
rect 34279 16836 34283 16892
rect 34283 16836 34339 16892
rect 34339 16836 34343 16892
rect 34279 16832 34343 16836
rect 34359 16892 34423 16896
rect 34359 16836 34363 16892
rect 34363 16836 34419 16892
rect 34419 16836 34423 16892
rect 34359 16832 34423 16836
rect 34439 16892 34503 16896
rect 34439 16836 34443 16892
rect 34443 16836 34499 16892
rect 34499 16836 34503 16892
rect 34439 16832 34503 16836
rect 34519 16892 34583 16896
rect 34519 16836 34523 16892
rect 34523 16836 34579 16892
rect 34579 16836 34583 16892
rect 34519 16832 34583 16836
rect 2820 16688 2884 16692
rect 2820 16632 2834 16688
rect 2834 16632 2884 16688
rect 2820 16628 2884 16632
rect 12204 16628 12268 16692
rect 19380 16628 19444 16692
rect 10474 16348 10538 16352
rect 10474 16292 10478 16348
rect 10478 16292 10534 16348
rect 10534 16292 10538 16348
rect 10474 16288 10538 16292
rect 10554 16348 10618 16352
rect 10554 16292 10558 16348
rect 10558 16292 10614 16348
rect 10614 16292 10618 16348
rect 10554 16288 10618 16292
rect 10634 16348 10698 16352
rect 10634 16292 10638 16348
rect 10638 16292 10694 16348
rect 10694 16292 10698 16348
rect 10634 16288 10698 16292
rect 10714 16348 10778 16352
rect 10714 16292 10718 16348
rect 10718 16292 10774 16348
rect 10774 16292 10778 16348
rect 10714 16288 10778 16292
rect 19996 16348 20060 16352
rect 19996 16292 20000 16348
rect 20000 16292 20056 16348
rect 20056 16292 20060 16348
rect 19996 16288 20060 16292
rect 20076 16348 20140 16352
rect 20076 16292 20080 16348
rect 20080 16292 20136 16348
rect 20136 16292 20140 16348
rect 20076 16288 20140 16292
rect 20156 16348 20220 16352
rect 20156 16292 20160 16348
rect 20160 16292 20216 16348
rect 20216 16292 20220 16348
rect 20156 16288 20220 16292
rect 20236 16348 20300 16352
rect 20236 16292 20240 16348
rect 20240 16292 20296 16348
rect 20296 16292 20300 16348
rect 20236 16288 20300 16292
rect 29518 16348 29582 16352
rect 29518 16292 29522 16348
rect 29522 16292 29578 16348
rect 29578 16292 29582 16348
rect 29518 16288 29582 16292
rect 29598 16348 29662 16352
rect 29598 16292 29602 16348
rect 29602 16292 29658 16348
rect 29658 16292 29662 16348
rect 29598 16288 29662 16292
rect 29678 16348 29742 16352
rect 29678 16292 29682 16348
rect 29682 16292 29738 16348
rect 29738 16292 29742 16348
rect 29678 16288 29742 16292
rect 29758 16348 29822 16352
rect 29758 16292 29762 16348
rect 29762 16292 29818 16348
rect 29818 16292 29822 16348
rect 29758 16288 29822 16292
rect 39040 16348 39104 16352
rect 39040 16292 39044 16348
rect 39044 16292 39100 16348
rect 39100 16292 39104 16348
rect 39040 16288 39104 16292
rect 39120 16348 39184 16352
rect 39120 16292 39124 16348
rect 39124 16292 39180 16348
rect 39180 16292 39184 16348
rect 39120 16288 39184 16292
rect 39200 16348 39264 16352
rect 39200 16292 39204 16348
rect 39204 16292 39260 16348
rect 39260 16292 39264 16348
rect 39200 16288 39264 16292
rect 39280 16348 39344 16352
rect 39280 16292 39284 16348
rect 39284 16292 39340 16348
rect 39340 16292 39344 16348
rect 39280 16288 39344 16292
rect 5713 15804 5777 15808
rect 5713 15748 5717 15804
rect 5717 15748 5773 15804
rect 5773 15748 5777 15804
rect 5713 15744 5777 15748
rect 5793 15804 5857 15808
rect 5793 15748 5797 15804
rect 5797 15748 5853 15804
rect 5853 15748 5857 15804
rect 5793 15744 5857 15748
rect 5873 15804 5937 15808
rect 5873 15748 5877 15804
rect 5877 15748 5933 15804
rect 5933 15748 5937 15804
rect 5873 15744 5937 15748
rect 5953 15804 6017 15808
rect 5953 15748 5957 15804
rect 5957 15748 6013 15804
rect 6013 15748 6017 15804
rect 5953 15744 6017 15748
rect 15235 15804 15299 15808
rect 15235 15748 15239 15804
rect 15239 15748 15295 15804
rect 15295 15748 15299 15804
rect 15235 15744 15299 15748
rect 15315 15804 15379 15808
rect 15315 15748 15319 15804
rect 15319 15748 15375 15804
rect 15375 15748 15379 15804
rect 15315 15744 15379 15748
rect 15395 15804 15459 15808
rect 15395 15748 15399 15804
rect 15399 15748 15455 15804
rect 15455 15748 15459 15804
rect 15395 15744 15459 15748
rect 15475 15804 15539 15808
rect 15475 15748 15479 15804
rect 15479 15748 15535 15804
rect 15535 15748 15539 15804
rect 15475 15744 15539 15748
rect 24757 15804 24821 15808
rect 24757 15748 24761 15804
rect 24761 15748 24817 15804
rect 24817 15748 24821 15804
rect 24757 15744 24821 15748
rect 24837 15804 24901 15808
rect 24837 15748 24841 15804
rect 24841 15748 24897 15804
rect 24897 15748 24901 15804
rect 24837 15744 24901 15748
rect 24917 15804 24981 15808
rect 24917 15748 24921 15804
rect 24921 15748 24977 15804
rect 24977 15748 24981 15804
rect 24917 15744 24981 15748
rect 24997 15804 25061 15808
rect 24997 15748 25001 15804
rect 25001 15748 25057 15804
rect 25057 15748 25061 15804
rect 24997 15744 25061 15748
rect 34279 15804 34343 15808
rect 34279 15748 34283 15804
rect 34283 15748 34339 15804
rect 34339 15748 34343 15804
rect 34279 15744 34343 15748
rect 34359 15804 34423 15808
rect 34359 15748 34363 15804
rect 34363 15748 34419 15804
rect 34419 15748 34423 15804
rect 34359 15744 34423 15748
rect 34439 15804 34503 15808
rect 34439 15748 34443 15804
rect 34443 15748 34499 15804
rect 34499 15748 34503 15804
rect 34439 15744 34503 15748
rect 34519 15804 34583 15808
rect 34519 15748 34523 15804
rect 34523 15748 34579 15804
rect 34579 15748 34583 15804
rect 34519 15744 34583 15748
rect 3188 15268 3252 15332
rect 4108 15268 4172 15332
rect 10474 15260 10538 15264
rect 10474 15204 10478 15260
rect 10478 15204 10534 15260
rect 10534 15204 10538 15260
rect 10474 15200 10538 15204
rect 10554 15260 10618 15264
rect 10554 15204 10558 15260
rect 10558 15204 10614 15260
rect 10614 15204 10618 15260
rect 10554 15200 10618 15204
rect 10634 15260 10698 15264
rect 10634 15204 10638 15260
rect 10638 15204 10694 15260
rect 10694 15204 10698 15260
rect 10634 15200 10698 15204
rect 10714 15260 10778 15264
rect 10714 15204 10718 15260
rect 10718 15204 10774 15260
rect 10774 15204 10778 15260
rect 10714 15200 10778 15204
rect 19996 15260 20060 15264
rect 19996 15204 20000 15260
rect 20000 15204 20056 15260
rect 20056 15204 20060 15260
rect 19996 15200 20060 15204
rect 20076 15260 20140 15264
rect 20076 15204 20080 15260
rect 20080 15204 20136 15260
rect 20136 15204 20140 15260
rect 20076 15200 20140 15204
rect 20156 15260 20220 15264
rect 20156 15204 20160 15260
rect 20160 15204 20216 15260
rect 20216 15204 20220 15260
rect 20156 15200 20220 15204
rect 20236 15260 20300 15264
rect 20236 15204 20240 15260
rect 20240 15204 20296 15260
rect 20296 15204 20300 15260
rect 20236 15200 20300 15204
rect 29518 15260 29582 15264
rect 29518 15204 29522 15260
rect 29522 15204 29578 15260
rect 29578 15204 29582 15260
rect 29518 15200 29582 15204
rect 29598 15260 29662 15264
rect 29598 15204 29602 15260
rect 29602 15204 29658 15260
rect 29658 15204 29662 15260
rect 29598 15200 29662 15204
rect 29678 15260 29742 15264
rect 29678 15204 29682 15260
rect 29682 15204 29738 15260
rect 29738 15204 29742 15260
rect 29678 15200 29742 15204
rect 29758 15260 29822 15264
rect 29758 15204 29762 15260
rect 29762 15204 29818 15260
rect 29818 15204 29822 15260
rect 29758 15200 29822 15204
rect 39040 15260 39104 15264
rect 39040 15204 39044 15260
rect 39044 15204 39100 15260
rect 39100 15204 39104 15260
rect 39040 15200 39104 15204
rect 39120 15260 39184 15264
rect 39120 15204 39124 15260
rect 39124 15204 39180 15260
rect 39180 15204 39184 15260
rect 39120 15200 39184 15204
rect 39200 15260 39264 15264
rect 39200 15204 39204 15260
rect 39204 15204 39260 15260
rect 39260 15204 39264 15260
rect 39200 15200 39264 15204
rect 39280 15260 39344 15264
rect 39280 15204 39284 15260
rect 39284 15204 39340 15260
rect 39340 15204 39344 15260
rect 39280 15200 39344 15204
rect 16436 15132 16500 15196
rect 19380 15132 19444 15196
rect 27476 15132 27540 15196
rect 12940 14996 13004 15060
rect 19564 14996 19628 15060
rect 20668 14724 20732 14788
rect 5713 14716 5777 14720
rect 5713 14660 5717 14716
rect 5717 14660 5773 14716
rect 5773 14660 5777 14716
rect 5713 14656 5777 14660
rect 5793 14716 5857 14720
rect 5793 14660 5797 14716
rect 5797 14660 5853 14716
rect 5853 14660 5857 14716
rect 5793 14656 5857 14660
rect 5873 14716 5937 14720
rect 5873 14660 5877 14716
rect 5877 14660 5933 14716
rect 5933 14660 5937 14716
rect 5873 14656 5937 14660
rect 5953 14716 6017 14720
rect 5953 14660 5957 14716
rect 5957 14660 6013 14716
rect 6013 14660 6017 14716
rect 5953 14656 6017 14660
rect 15235 14716 15299 14720
rect 15235 14660 15239 14716
rect 15239 14660 15295 14716
rect 15295 14660 15299 14716
rect 15235 14656 15299 14660
rect 15315 14716 15379 14720
rect 15315 14660 15319 14716
rect 15319 14660 15375 14716
rect 15375 14660 15379 14716
rect 15315 14656 15379 14660
rect 15395 14716 15459 14720
rect 15395 14660 15399 14716
rect 15399 14660 15455 14716
rect 15455 14660 15459 14716
rect 15395 14656 15459 14660
rect 15475 14716 15539 14720
rect 15475 14660 15479 14716
rect 15479 14660 15535 14716
rect 15535 14660 15539 14716
rect 15475 14656 15539 14660
rect 24757 14716 24821 14720
rect 24757 14660 24761 14716
rect 24761 14660 24817 14716
rect 24817 14660 24821 14716
rect 24757 14656 24821 14660
rect 24837 14716 24901 14720
rect 24837 14660 24841 14716
rect 24841 14660 24897 14716
rect 24897 14660 24901 14716
rect 24837 14656 24901 14660
rect 24917 14716 24981 14720
rect 24917 14660 24921 14716
rect 24921 14660 24977 14716
rect 24977 14660 24981 14716
rect 24917 14656 24981 14660
rect 24997 14716 25061 14720
rect 24997 14660 25001 14716
rect 25001 14660 25057 14716
rect 25057 14660 25061 14716
rect 24997 14656 25061 14660
rect 34279 14716 34343 14720
rect 34279 14660 34283 14716
rect 34283 14660 34339 14716
rect 34339 14660 34343 14716
rect 34279 14656 34343 14660
rect 34359 14716 34423 14720
rect 34359 14660 34363 14716
rect 34363 14660 34419 14716
rect 34419 14660 34423 14716
rect 34359 14656 34423 14660
rect 34439 14716 34503 14720
rect 34439 14660 34443 14716
rect 34443 14660 34499 14716
rect 34499 14660 34503 14716
rect 34439 14656 34503 14660
rect 34519 14716 34583 14720
rect 34519 14660 34523 14716
rect 34523 14660 34579 14716
rect 34579 14660 34583 14716
rect 34519 14656 34583 14660
rect 10474 14172 10538 14176
rect 10474 14116 10478 14172
rect 10478 14116 10534 14172
rect 10534 14116 10538 14172
rect 10474 14112 10538 14116
rect 10554 14172 10618 14176
rect 10554 14116 10558 14172
rect 10558 14116 10614 14172
rect 10614 14116 10618 14172
rect 10554 14112 10618 14116
rect 10634 14172 10698 14176
rect 10634 14116 10638 14172
rect 10638 14116 10694 14172
rect 10694 14116 10698 14172
rect 10634 14112 10698 14116
rect 10714 14172 10778 14176
rect 10714 14116 10718 14172
rect 10718 14116 10774 14172
rect 10774 14116 10778 14172
rect 10714 14112 10778 14116
rect 19996 14172 20060 14176
rect 19996 14116 20000 14172
rect 20000 14116 20056 14172
rect 20056 14116 20060 14172
rect 19996 14112 20060 14116
rect 20076 14172 20140 14176
rect 20076 14116 20080 14172
rect 20080 14116 20136 14172
rect 20136 14116 20140 14172
rect 20076 14112 20140 14116
rect 20156 14172 20220 14176
rect 20156 14116 20160 14172
rect 20160 14116 20216 14172
rect 20216 14116 20220 14172
rect 20156 14112 20220 14116
rect 20236 14172 20300 14176
rect 20236 14116 20240 14172
rect 20240 14116 20296 14172
rect 20296 14116 20300 14172
rect 20236 14112 20300 14116
rect 29518 14172 29582 14176
rect 29518 14116 29522 14172
rect 29522 14116 29578 14172
rect 29578 14116 29582 14172
rect 29518 14112 29582 14116
rect 29598 14172 29662 14176
rect 29598 14116 29602 14172
rect 29602 14116 29658 14172
rect 29658 14116 29662 14172
rect 29598 14112 29662 14116
rect 29678 14172 29742 14176
rect 29678 14116 29682 14172
rect 29682 14116 29738 14172
rect 29738 14116 29742 14172
rect 29678 14112 29742 14116
rect 29758 14172 29822 14176
rect 29758 14116 29762 14172
rect 29762 14116 29818 14172
rect 29818 14116 29822 14172
rect 29758 14112 29822 14116
rect 39040 14172 39104 14176
rect 39040 14116 39044 14172
rect 39044 14116 39100 14172
rect 39100 14116 39104 14172
rect 39040 14112 39104 14116
rect 39120 14172 39184 14176
rect 39120 14116 39124 14172
rect 39124 14116 39180 14172
rect 39180 14116 39184 14172
rect 39120 14112 39184 14116
rect 39200 14172 39264 14176
rect 39200 14116 39204 14172
rect 39204 14116 39260 14172
rect 39260 14116 39264 14172
rect 39200 14112 39264 14116
rect 39280 14172 39344 14176
rect 39280 14116 39284 14172
rect 39284 14116 39340 14172
rect 39340 14116 39344 14172
rect 39280 14112 39344 14116
rect 12572 13908 12636 13972
rect 14596 13908 14660 13972
rect 16804 13636 16868 13700
rect 5713 13628 5777 13632
rect 5713 13572 5717 13628
rect 5717 13572 5773 13628
rect 5773 13572 5777 13628
rect 5713 13568 5777 13572
rect 5793 13628 5857 13632
rect 5793 13572 5797 13628
rect 5797 13572 5853 13628
rect 5853 13572 5857 13628
rect 5793 13568 5857 13572
rect 5873 13628 5937 13632
rect 5873 13572 5877 13628
rect 5877 13572 5933 13628
rect 5933 13572 5937 13628
rect 5873 13568 5937 13572
rect 5953 13628 6017 13632
rect 5953 13572 5957 13628
rect 5957 13572 6013 13628
rect 6013 13572 6017 13628
rect 5953 13568 6017 13572
rect 15235 13628 15299 13632
rect 15235 13572 15239 13628
rect 15239 13572 15295 13628
rect 15295 13572 15299 13628
rect 15235 13568 15299 13572
rect 15315 13628 15379 13632
rect 15315 13572 15319 13628
rect 15319 13572 15375 13628
rect 15375 13572 15379 13628
rect 15315 13568 15379 13572
rect 15395 13628 15459 13632
rect 15395 13572 15399 13628
rect 15399 13572 15455 13628
rect 15455 13572 15459 13628
rect 15395 13568 15459 13572
rect 15475 13628 15539 13632
rect 15475 13572 15479 13628
rect 15479 13572 15535 13628
rect 15535 13572 15539 13628
rect 15475 13568 15539 13572
rect 24757 13628 24821 13632
rect 24757 13572 24761 13628
rect 24761 13572 24817 13628
rect 24817 13572 24821 13628
rect 24757 13568 24821 13572
rect 24837 13628 24901 13632
rect 24837 13572 24841 13628
rect 24841 13572 24897 13628
rect 24897 13572 24901 13628
rect 24837 13568 24901 13572
rect 24917 13628 24981 13632
rect 24917 13572 24921 13628
rect 24921 13572 24977 13628
rect 24977 13572 24981 13628
rect 24917 13568 24981 13572
rect 24997 13628 25061 13632
rect 24997 13572 25001 13628
rect 25001 13572 25057 13628
rect 25057 13572 25061 13628
rect 24997 13568 25061 13572
rect 34279 13628 34343 13632
rect 34279 13572 34283 13628
rect 34283 13572 34339 13628
rect 34339 13572 34343 13628
rect 34279 13568 34343 13572
rect 34359 13628 34423 13632
rect 34359 13572 34363 13628
rect 34363 13572 34419 13628
rect 34419 13572 34423 13628
rect 34359 13568 34423 13572
rect 34439 13628 34503 13632
rect 34439 13572 34443 13628
rect 34443 13572 34499 13628
rect 34499 13572 34503 13628
rect 34439 13568 34503 13572
rect 34519 13628 34583 13632
rect 34519 13572 34523 13628
rect 34523 13572 34579 13628
rect 34579 13572 34583 13628
rect 34519 13568 34583 13572
rect 14780 13500 14844 13564
rect 15700 13500 15764 13564
rect 18828 13560 18892 13564
rect 18828 13504 18842 13560
rect 18842 13504 18892 13560
rect 18828 13500 18892 13504
rect 28396 13500 28460 13564
rect 30420 13500 30484 13564
rect 27844 13228 27908 13292
rect 30052 13228 30116 13292
rect 10474 13084 10538 13088
rect 10474 13028 10478 13084
rect 10478 13028 10534 13084
rect 10534 13028 10538 13084
rect 10474 13024 10538 13028
rect 10554 13084 10618 13088
rect 10554 13028 10558 13084
rect 10558 13028 10614 13084
rect 10614 13028 10618 13084
rect 10554 13024 10618 13028
rect 10634 13084 10698 13088
rect 10634 13028 10638 13084
rect 10638 13028 10694 13084
rect 10694 13028 10698 13084
rect 10634 13024 10698 13028
rect 10714 13084 10778 13088
rect 10714 13028 10718 13084
rect 10718 13028 10774 13084
rect 10774 13028 10778 13084
rect 10714 13024 10778 13028
rect 19996 13084 20060 13088
rect 19996 13028 20000 13084
rect 20000 13028 20056 13084
rect 20056 13028 20060 13084
rect 19996 13024 20060 13028
rect 20076 13084 20140 13088
rect 20076 13028 20080 13084
rect 20080 13028 20136 13084
rect 20136 13028 20140 13084
rect 20076 13024 20140 13028
rect 20156 13084 20220 13088
rect 20156 13028 20160 13084
rect 20160 13028 20216 13084
rect 20216 13028 20220 13084
rect 20156 13024 20220 13028
rect 20236 13084 20300 13088
rect 20236 13028 20240 13084
rect 20240 13028 20296 13084
rect 20296 13028 20300 13084
rect 20236 13024 20300 13028
rect 29518 13084 29582 13088
rect 29518 13028 29522 13084
rect 29522 13028 29578 13084
rect 29578 13028 29582 13084
rect 29518 13024 29582 13028
rect 29598 13084 29662 13088
rect 29598 13028 29602 13084
rect 29602 13028 29658 13084
rect 29658 13028 29662 13084
rect 29598 13024 29662 13028
rect 29678 13084 29742 13088
rect 29678 13028 29682 13084
rect 29682 13028 29738 13084
rect 29738 13028 29742 13084
rect 29678 13024 29742 13028
rect 29758 13084 29822 13088
rect 29758 13028 29762 13084
rect 29762 13028 29818 13084
rect 29818 13028 29822 13084
rect 29758 13024 29822 13028
rect 39040 13084 39104 13088
rect 39040 13028 39044 13084
rect 39044 13028 39100 13084
rect 39100 13028 39104 13084
rect 39040 13024 39104 13028
rect 39120 13084 39184 13088
rect 39120 13028 39124 13084
rect 39124 13028 39180 13084
rect 39180 13028 39184 13084
rect 39120 13024 39184 13028
rect 39200 13084 39264 13088
rect 39200 13028 39204 13084
rect 39204 13028 39260 13084
rect 39260 13028 39264 13084
rect 39200 13024 39264 13028
rect 39280 13084 39344 13088
rect 39280 13028 39284 13084
rect 39284 13028 39340 13084
rect 39340 13028 39344 13084
rect 39280 13024 39344 13028
rect 15700 12956 15764 13020
rect 8892 12684 8956 12748
rect 5396 12548 5460 12612
rect 19564 12684 19628 12748
rect 15700 12548 15764 12612
rect 5713 12540 5777 12544
rect 5713 12484 5717 12540
rect 5717 12484 5773 12540
rect 5773 12484 5777 12540
rect 5713 12480 5777 12484
rect 5793 12540 5857 12544
rect 5793 12484 5797 12540
rect 5797 12484 5853 12540
rect 5853 12484 5857 12540
rect 5793 12480 5857 12484
rect 5873 12540 5937 12544
rect 5873 12484 5877 12540
rect 5877 12484 5933 12540
rect 5933 12484 5937 12540
rect 5873 12480 5937 12484
rect 5953 12540 6017 12544
rect 5953 12484 5957 12540
rect 5957 12484 6013 12540
rect 6013 12484 6017 12540
rect 5953 12480 6017 12484
rect 15235 12540 15299 12544
rect 15235 12484 15239 12540
rect 15239 12484 15295 12540
rect 15295 12484 15299 12540
rect 15235 12480 15299 12484
rect 15315 12540 15379 12544
rect 15315 12484 15319 12540
rect 15319 12484 15375 12540
rect 15375 12484 15379 12540
rect 15315 12480 15379 12484
rect 15395 12540 15459 12544
rect 15395 12484 15399 12540
rect 15399 12484 15455 12540
rect 15455 12484 15459 12540
rect 15395 12480 15459 12484
rect 15475 12540 15539 12544
rect 15475 12484 15479 12540
rect 15479 12484 15535 12540
rect 15535 12484 15539 12540
rect 15475 12480 15539 12484
rect 24757 12540 24821 12544
rect 24757 12484 24761 12540
rect 24761 12484 24817 12540
rect 24817 12484 24821 12540
rect 24757 12480 24821 12484
rect 24837 12540 24901 12544
rect 24837 12484 24841 12540
rect 24841 12484 24897 12540
rect 24897 12484 24901 12540
rect 24837 12480 24901 12484
rect 24917 12540 24981 12544
rect 24917 12484 24921 12540
rect 24921 12484 24977 12540
rect 24977 12484 24981 12540
rect 24917 12480 24981 12484
rect 24997 12540 25061 12544
rect 24997 12484 25001 12540
rect 25001 12484 25057 12540
rect 25057 12484 25061 12540
rect 24997 12480 25061 12484
rect 34279 12540 34343 12544
rect 34279 12484 34283 12540
rect 34283 12484 34339 12540
rect 34339 12484 34343 12540
rect 34279 12480 34343 12484
rect 34359 12540 34423 12544
rect 34359 12484 34363 12540
rect 34363 12484 34419 12540
rect 34419 12484 34423 12540
rect 34359 12480 34423 12484
rect 34439 12540 34503 12544
rect 34439 12484 34443 12540
rect 34443 12484 34499 12540
rect 34499 12484 34503 12540
rect 34439 12480 34503 12484
rect 34519 12540 34583 12544
rect 34519 12484 34523 12540
rect 34523 12484 34579 12540
rect 34579 12484 34583 12540
rect 34519 12480 34583 12484
rect 31708 12412 31772 12476
rect 14596 12276 14660 12340
rect 16436 12276 16500 12340
rect 23428 12140 23492 12204
rect 31156 12140 31220 12204
rect 9444 12064 9508 12068
rect 9444 12008 9458 12064
rect 9458 12008 9508 12064
rect 9444 12004 9508 12008
rect 13860 12004 13924 12068
rect 17724 12004 17788 12068
rect 10474 11996 10538 12000
rect 10474 11940 10478 11996
rect 10478 11940 10534 11996
rect 10534 11940 10538 11996
rect 10474 11936 10538 11940
rect 10554 11996 10618 12000
rect 10554 11940 10558 11996
rect 10558 11940 10614 11996
rect 10614 11940 10618 11996
rect 10554 11936 10618 11940
rect 10634 11996 10698 12000
rect 10634 11940 10638 11996
rect 10638 11940 10694 11996
rect 10694 11940 10698 11996
rect 10634 11936 10698 11940
rect 10714 11996 10778 12000
rect 10714 11940 10718 11996
rect 10718 11940 10774 11996
rect 10774 11940 10778 11996
rect 10714 11936 10778 11940
rect 19996 11996 20060 12000
rect 19996 11940 20000 11996
rect 20000 11940 20056 11996
rect 20056 11940 20060 11996
rect 19996 11936 20060 11940
rect 20076 11996 20140 12000
rect 20076 11940 20080 11996
rect 20080 11940 20136 11996
rect 20136 11940 20140 11996
rect 20076 11936 20140 11940
rect 20156 11996 20220 12000
rect 20156 11940 20160 11996
rect 20160 11940 20216 11996
rect 20216 11940 20220 11996
rect 20156 11936 20220 11940
rect 20236 11996 20300 12000
rect 20236 11940 20240 11996
rect 20240 11940 20296 11996
rect 20296 11940 20300 11996
rect 20236 11936 20300 11940
rect 9628 11868 9692 11932
rect 25820 11792 25884 11796
rect 25820 11736 25834 11792
rect 25834 11736 25884 11792
rect 25820 11732 25884 11736
rect 26740 11732 26804 11796
rect 29518 11996 29582 12000
rect 29518 11940 29522 11996
rect 29522 11940 29578 11996
rect 29578 11940 29582 11996
rect 29518 11936 29582 11940
rect 29598 11996 29662 12000
rect 29598 11940 29602 11996
rect 29602 11940 29658 11996
rect 29658 11940 29662 11996
rect 29598 11936 29662 11940
rect 29678 11996 29742 12000
rect 29678 11940 29682 11996
rect 29682 11940 29738 11996
rect 29738 11940 29742 11996
rect 29678 11936 29742 11940
rect 29758 11996 29822 12000
rect 29758 11940 29762 11996
rect 29762 11940 29818 11996
rect 29818 11940 29822 11996
rect 29758 11936 29822 11940
rect 39040 11996 39104 12000
rect 39040 11940 39044 11996
rect 39044 11940 39100 11996
rect 39100 11940 39104 11996
rect 39040 11936 39104 11940
rect 39120 11996 39184 12000
rect 39120 11940 39124 11996
rect 39124 11940 39180 11996
rect 39180 11940 39184 11996
rect 39120 11936 39184 11940
rect 39200 11996 39264 12000
rect 39200 11940 39204 11996
rect 39204 11940 39260 11996
rect 39260 11940 39264 11996
rect 39200 11936 39264 11940
rect 39280 11996 39344 12000
rect 39280 11940 39284 11996
rect 39284 11940 39340 11996
rect 39340 11940 39344 11996
rect 39280 11936 39344 11940
rect 28212 11596 28276 11660
rect 11100 11460 11164 11524
rect 5713 11452 5777 11456
rect 5713 11396 5717 11452
rect 5717 11396 5773 11452
rect 5773 11396 5777 11452
rect 5713 11392 5777 11396
rect 5793 11452 5857 11456
rect 5793 11396 5797 11452
rect 5797 11396 5853 11452
rect 5853 11396 5857 11452
rect 5793 11392 5857 11396
rect 5873 11452 5937 11456
rect 5873 11396 5877 11452
rect 5877 11396 5933 11452
rect 5933 11396 5937 11452
rect 5873 11392 5937 11396
rect 5953 11452 6017 11456
rect 5953 11396 5957 11452
rect 5957 11396 6013 11452
rect 6013 11396 6017 11452
rect 5953 11392 6017 11396
rect 15235 11452 15299 11456
rect 15235 11396 15239 11452
rect 15239 11396 15295 11452
rect 15295 11396 15299 11452
rect 15235 11392 15299 11396
rect 15315 11452 15379 11456
rect 15315 11396 15319 11452
rect 15319 11396 15375 11452
rect 15375 11396 15379 11452
rect 15315 11392 15379 11396
rect 15395 11452 15459 11456
rect 15395 11396 15399 11452
rect 15399 11396 15455 11452
rect 15455 11396 15459 11452
rect 15395 11392 15459 11396
rect 15475 11452 15539 11456
rect 15475 11396 15479 11452
rect 15479 11396 15535 11452
rect 15535 11396 15539 11452
rect 15475 11392 15539 11396
rect 24757 11452 24821 11456
rect 24757 11396 24761 11452
rect 24761 11396 24817 11452
rect 24817 11396 24821 11452
rect 24757 11392 24821 11396
rect 24837 11452 24901 11456
rect 24837 11396 24841 11452
rect 24841 11396 24897 11452
rect 24897 11396 24901 11452
rect 24837 11392 24901 11396
rect 24917 11452 24981 11456
rect 24917 11396 24921 11452
rect 24921 11396 24977 11452
rect 24977 11396 24981 11452
rect 24917 11392 24981 11396
rect 24997 11452 25061 11456
rect 24997 11396 25001 11452
rect 25001 11396 25057 11452
rect 25057 11396 25061 11452
rect 24997 11392 25061 11396
rect 34279 11452 34343 11456
rect 34279 11396 34283 11452
rect 34283 11396 34339 11452
rect 34339 11396 34343 11452
rect 34279 11392 34343 11396
rect 34359 11452 34423 11456
rect 34359 11396 34363 11452
rect 34363 11396 34419 11452
rect 34419 11396 34423 11452
rect 34359 11392 34423 11396
rect 34439 11452 34503 11456
rect 34439 11396 34443 11452
rect 34443 11396 34499 11452
rect 34499 11396 34503 11452
rect 34439 11392 34503 11396
rect 34519 11452 34583 11456
rect 34519 11396 34523 11452
rect 34523 11396 34579 11452
rect 34579 11396 34583 11452
rect 34519 11392 34583 11396
rect 9812 11324 9876 11388
rect 7604 11188 7668 11252
rect 9996 11188 10060 11252
rect 10180 11112 10244 11116
rect 10180 11056 10230 11112
rect 10230 11056 10244 11112
rect 10180 11052 10244 11056
rect 10474 10908 10538 10912
rect 10474 10852 10478 10908
rect 10478 10852 10534 10908
rect 10534 10852 10538 10908
rect 10474 10848 10538 10852
rect 10554 10908 10618 10912
rect 10554 10852 10558 10908
rect 10558 10852 10614 10908
rect 10614 10852 10618 10908
rect 10554 10848 10618 10852
rect 10634 10908 10698 10912
rect 10634 10852 10638 10908
rect 10638 10852 10694 10908
rect 10694 10852 10698 10908
rect 10634 10848 10698 10852
rect 10714 10908 10778 10912
rect 10714 10852 10718 10908
rect 10718 10852 10774 10908
rect 10774 10852 10778 10908
rect 10714 10848 10778 10852
rect 12020 10976 12084 10980
rect 12020 10920 12070 10976
rect 12070 10920 12084 10976
rect 12020 10916 12084 10920
rect 16068 11052 16132 11116
rect 16804 11052 16868 11116
rect 16988 11112 17052 11116
rect 16988 11056 17002 11112
rect 17002 11056 17052 11112
rect 16988 11052 17052 11056
rect 31156 11112 31220 11116
rect 31156 11056 31206 11112
rect 31206 11056 31220 11112
rect 31156 11052 31220 11056
rect 12940 10780 13004 10844
rect 14412 10840 14476 10844
rect 14412 10784 14462 10840
rect 14462 10784 14476 10840
rect 14412 10780 14476 10784
rect 15700 10780 15764 10844
rect 25452 10916 25516 10980
rect 19996 10908 20060 10912
rect 19996 10852 20000 10908
rect 20000 10852 20056 10908
rect 20056 10852 20060 10908
rect 19996 10848 20060 10852
rect 20076 10908 20140 10912
rect 20076 10852 20080 10908
rect 20080 10852 20136 10908
rect 20136 10852 20140 10908
rect 20076 10848 20140 10852
rect 20156 10908 20220 10912
rect 20156 10852 20160 10908
rect 20160 10852 20216 10908
rect 20216 10852 20220 10908
rect 20156 10848 20220 10852
rect 20236 10908 20300 10912
rect 20236 10852 20240 10908
rect 20240 10852 20296 10908
rect 20296 10852 20300 10908
rect 20236 10848 20300 10852
rect 29316 10916 29380 10980
rect 29518 10908 29582 10912
rect 29518 10852 29522 10908
rect 29522 10852 29578 10908
rect 29578 10852 29582 10908
rect 29518 10848 29582 10852
rect 29598 10908 29662 10912
rect 29598 10852 29602 10908
rect 29602 10852 29658 10908
rect 29658 10852 29662 10908
rect 29598 10848 29662 10852
rect 29678 10908 29742 10912
rect 29678 10852 29682 10908
rect 29682 10852 29738 10908
rect 29738 10852 29742 10908
rect 29678 10848 29742 10852
rect 29758 10908 29822 10912
rect 29758 10852 29762 10908
rect 29762 10852 29818 10908
rect 29818 10852 29822 10908
rect 29758 10848 29822 10852
rect 39040 10908 39104 10912
rect 39040 10852 39044 10908
rect 39044 10852 39100 10908
rect 39100 10852 39104 10908
rect 39040 10848 39104 10852
rect 39120 10908 39184 10912
rect 39120 10852 39124 10908
rect 39124 10852 39180 10908
rect 39180 10852 39184 10908
rect 39120 10848 39184 10852
rect 39200 10908 39264 10912
rect 39200 10852 39204 10908
rect 39204 10852 39260 10908
rect 39260 10852 39264 10908
rect 39200 10848 39264 10852
rect 39280 10908 39344 10912
rect 39280 10852 39284 10908
rect 39284 10852 39340 10908
rect 39340 10852 39344 10908
rect 39280 10848 39344 10852
rect 27476 10840 27540 10844
rect 27476 10784 27526 10840
rect 27526 10784 27540 10840
rect 27476 10780 27540 10784
rect 29316 10508 29380 10572
rect 5713 10364 5777 10368
rect 5713 10308 5717 10364
rect 5717 10308 5773 10364
rect 5773 10308 5777 10364
rect 5713 10304 5777 10308
rect 5793 10364 5857 10368
rect 5793 10308 5797 10364
rect 5797 10308 5853 10364
rect 5853 10308 5857 10364
rect 5793 10304 5857 10308
rect 5873 10364 5937 10368
rect 5873 10308 5877 10364
rect 5877 10308 5933 10364
rect 5933 10308 5937 10364
rect 5873 10304 5937 10308
rect 5953 10364 6017 10368
rect 5953 10308 5957 10364
rect 5957 10308 6013 10364
rect 6013 10308 6017 10364
rect 5953 10304 6017 10308
rect 15235 10364 15299 10368
rect 15235 10308 15239 10364
rect 15239 10308 15295 10364
rect 15295 10308 15299 10364
rect 15235 10304 15299 10308
rect 15315 10364 15379 10368
rect 15315 10308 15319 10364
rect 15319 10308 15375 10364
rect 15375 10308 15379 10364
rect 15315 10304 15379 10308
rect 15395 10364 15459 10368
rect 15395 10308 15399 10364
rect 15399 10308 15455 10364
rect 15455 10308 15459 10364
rect 15395 10304 15459 10308
rect 15475 10364 15539 10368
rect 15475 10308 15479 10364
rect 15479 10308 15535 10364
rect 15535 10308 15539 10364
rect 15475 10304 15539 10308
rect 24757 10364 24821 10368
rect 24757 10308 24761 10364
rect 24761 10308 24817 10364
rect 24817 10308 24821 10364
rect 24757 10304 24821 10308
rect 24837 10364 24901 10368
rect 24837 10308 24841 10364
rect 24841 10308 24897 10364
rect 24897 10308 24901 10364
rect 24837 10304 24901 10308
rect 24917 10364 24981 10368
rect 24917 10308 24921 10364
rect 24921 10308 24977 10364
rect 24977 10308 24981 10364
rect 24917 10304 24981 10308
rect 24997 10364 25061 10368
rect 24997 10308 25001 10364
rect 25001 10308 25057 10364
rect 25057 10308 25061 10364
rect 24997 10304 25061 10308
rect 34279 10364 34343 10368
rect 34279 10308 34283 10364
rect 34283 10308 34339 10364
rect 34339 10308 34343 10364
rect 34279 10304 34343 10308
rect 34359 10364 34423 10368
rect 34359 10308 34363 10364
rect 34363 10308 34419 10364
rect 34419 10308 34423 10364
rect 34359 10304 34423 10308
rect 34439 10364 34503 10368
rect 34439 10308 34443 10364
rect 34443 10308 34499 10364
rect 34499 10308 34503 10364
rect 34439 10304 34503 10308
rect 34519 10364 34583 10368
rect 34519 10308 34523 10364
rect 34523 10308 34579 10364
rect 34579 10308 34583 10364
rect 34519 10304 34583 10308
rect 28948 10100 29012 10164
rect 9812 9888 9876 9892
rect 9812 9832 9826 9888
rect 9826 9832 9876 9888
rect 9812 9828 9876 9832
rect 12020 9888 12084 9892
rect 12020 9832 12070 9888
rect 12070 9832 12084 9888
rect 12020 9828 12084 9832
rect 10474 9820 10538 9824
rect 10474 9764 10478 9820
rect 10478 9764 10534 9820
rect 10534 9764 10538 9820
rect 10474 9760 10538 9764
rect 10554 9820 10618 9824
rect 10554 9764 10558 9820
rect 10558 9764 10614 9820
rect 10614 9764 10618 9820
rect 10554 9760 10618 9764
rect 10634 9820 10698 9824
rect 10634 9764 10638 9820
rect 10638 9764 10694 9820
rect 10694 9764 10698 9820
rect 10634 9760 10698 9764
rect 10714 9820 10778 9824
rect 10714 9764 10718 9820
rect 10718 9764 10774 9820
rect 10774 9764 10778 9820
rect 10714 9760 10778 9764
rect 2636 9752 2700 9756
rect 2636 9696 2650 9752
rect 2650 9696 2700 9752
rect 2636 9692 2700 9696
rect 9996 9692 10060 9756
rect 29132 9828 29196 9892
rect 19996 9820 20060 9824
rect 19996 9764 20000 9820
rect 20000 9764 20056 9820
rect 20056 9764 20060 9820
rect 19996 9760 20060 9764
rect 20076 9820 20140 9824
rect 20076 9764 20080 9820
rect 20080 9764 20136 9820
rect 20136 9764 20140 9820
rect 20076 9760 20140 9764
rect 20156 9820 20220 9824
rect 20156 9764 20160 9820
rect 20160 9764 20216 9820
rect 20216 9764 20220 9820
rect 20156 9760 20220 9764
rect 20236 9820 20300 9824
rect 20236 9764 20240 9820
rect 20240 9764 20296 9820
rect 20296 9764 20300 9820
rect 20236 9760 20300 9764
rect 29518 9820 29582 9824
rect 29518 9764 29522 9820
rect 29522 9764 29578 9820
rect 29578 9764 29582 9820
rect 29518 9760 29582 9764
rect 29598 9820 29662 9824
rect 29598 9764 29602 9820
rect 29602 9764 29658 9820
rect 29658 9764 29662 9820
rect 29598 9760 29662 9764
rect 29678 9820 29742 9824
rect 29678 9764 29682 9820
rect 29682 9764 29738 9820
rect 29738 9764 29742 9820
rect 29678 9760 29742 9764
rect 29758 9820 29822 9824
rect 29758 9764 29762 9820
rect 29762 9764 29818 9820
rect 29818 9764 29822 9820
rect 29758 9760 29822 9764
rect 39040 9820 39104 9824
rect 39040 9764 39044 9820
rect 39044 9764 39100 9820
rect 39100 9764 39104 9820
rect 39040 9760 39104 9764
rect 39120 9820 39184 9824
rect 39120 9764 39124 9820
rect 39124 9764 39180 9820
rect 39180 9764 39184 9820
rect 39120 9760 39184 9764
rect 39200 9820 39264 9824
rect 39200 9764 39204 9820
rect 39204 9764 39260 9820
rect 39260 9764 39264 9820
rect 39200 9760 39264 9764
rect 39280 9820 39344 9824
rect 39280 9764 39284 9820
rect 39284 9764 39340 9820
rect 39340 9764 39344 9820
rect 39280 9760 39344 9764
rect 12756 9556 12820 9620
rect 13124 9556 13188 9620
rect 15700 9556 15764 9620
rect 26924 9692 26988 9756
rect 27844 9752 27908 9756
rect 27844 9696 27894 9752
rect 27894 9696 27908 9752
rect 27844 9692 27908 9696
rect 30236 9752 30300 9756
rect 30236 9696 30250 9752
rect 30250 9696 30300 9752
rect 22692 9616 22756 9620
rect 22692 9560 22742 9616
rect 22742 9560 22756 9616
rect 22692 9556 22756 9560
rect 28580 9556 28644 9620
rect 30236 9692 30300 9696
rect 31340 9752 31404 9756
rect 31340 9696 31390 9752
rect 31390 9696 31404 9752
rect 31340 9692 31404 9696
rect 31892 9556 31956 9620
rect 13492 9420 13556 9484
rect 14044 9284 14108 9348
rect 27844 9420 27908 9484
rect 28028 9420 28092 9484
rect 28764 9284 28828 9348
rect 5713 9276 5777 9280
rect 5713 9220 5717 9276
rect 5717 9220 5773 9276
rect 5773 9220 5777 9276
rect 5713 9216 5777 9220
rect 5793 9276 5857 9280
rect 5793 9220 5797 9276
rect 5797 9220 5853 9276
rect 5853 9220 5857 9276
rect 5793 9216 5857 9220
rect 5873 9276 5937 9280
rect 5873 9220 5877 9276
rect 5877 9220 5933 9276
rect 5933 9220 5937 9276
rect 5873 9216 5937 9220
rect 5953 9276 6017 9280
rect 5953 9220 5957 9276
rect 5957 9220 6013 9276
rect 6013 9220 6017 9276
rect 5953 9216 6017 9220
rect 15235 9276 15299 9280
rect 15235 9220 15239 9276
rect 15239 9220 15295 9276
rect 15295 9220 15299 9276
rect 15235 9216 15299 9220
rect 15315 9276 15379 9280
rect 15315 9220 15319 9276
rect 15319 9220 15375 9276
rect 15375 9220 15379 9276
rect 15315 9216 15379 9220
rect 15395 9276 15459 9280
rect 15395 9220 15399 9276
rect 15399 9220 15455 9276
rect 15455 9220 15459 9276
rect 15395 9216 15459 9220
rect 15475 9276 15539 9280
rect 15475 9220 15479 9276
rect 15479 9220 15535 9276
rect 15535 9220 15539 9276
rect 15475 9216 15539 9220
rect 24757 9276 24821 9280
rect 24757 9220 24761 9276
rect 24761 9220 24817 9276
rect 24817 9220 24821 9276
rect 24757 9216 24821 9220
rect 24837 9276 24901 9280
rect 24837 9220 24841 9276
rect 24841 9220 24897 9276
rect 24897 9220 24901 9276
rect 24837 9216 24901 9220
rect 24917 9276 24981 9280
rect 24917 9220 24921 9276
rect 24921 9220 24977 9276
rect 24977 9220 24981 9276
rect 24917 9216 24981 9220
rect 24997 9276 25061 9280
rect 24997 9220 25001 9276
rect 25001 9220 25057 9276
rect 25057 9220 25061 9276
rect 24997 9216 25061 9220
rect 34279 9276 34343 9280
rect 34279 9220 34283 9276
rect 34283 9220 34339 9276
rect 34339 9220 34343 9276
rect 34279 9216 34343 9220
rect 34359 9276 34423 9280
rect 34359 9220 34363 9276
rect 34363 9220 34419 9276
rect 34419 9220 34423 9276
rect 34359 9216 34423 9220
rect 34439 9276 34503 9280
rect 34439 9220 34443 9276
rect 34443 9220 34499 9276
rect 34499 9220 34503 9276
rect 34439 9216 34503 9220
rect 34519 9276 34583 9280
rect 34519 9220 34523 9276
rect 34523 9220 34579 9276
rect 34579 9220 34583 9276
rect 34519 9216 34583 9220
rect 15102 9072 15166 9076
rect 15102 9016 15106 9072
rect 15106 9016 15162 9072
rect 15162 9016 15166 9072
rect 15102 9012 15166 9016
rect 30420 9148 30484 9212
rect 18644 8876 18708 8940
rect 20668 8740 20732 8804
rect 24532 8876 24596 8940
rect 34652 8876 34716 8940
rect 28764 8740 28828 8804
rect 32812 8740 32876 8804
rect 32996 8740 33060 8804
rect 10474 8732 10538 8736
rect 10474 8676 10478 8732
rect 10478 8676 10534 8732
rect 10534 8676 10538 8732
rect 10474 8672 10538 8676
rect 10554 8732 10618 8736
rect 10554 8676 10558 8732
rect 10558 8676 10614 8732
rect 10614 8676 10618 8732
rect 10554 8672 10618 8676
rect 10634 8732 10698 8736
rect 10634 8676 10638 8732
rect 10638 8676 10694 8732
rect 10694 8676 10698 8732
rect 10634 8672 10698 8676
rect 10714 8732 10778 8736
rect 10714 8676 10718 8732
rect 10718 8676 10774 8732
rect 10774 8676 10778 8732
rect 10714 8672 10778 8676
rect 19996 8732 20060 8736
rect 19996 8676 20000 8732
rect 20000 8676 20056 8732
rect 20056 8676 20060 8732
rect 19996 8672 20060 8676
rect 20076 8732 20140 8736
rect 20076 8676 20080 8732
rect 20080 8676 20136 8732
rect 20136 8676 20140 8732
rect 20076 8672 20140 8676
rect 20156 8732 20220 8736
rect 20156 8676 20160 8732
rect 20160 8676 20216 8732
rect 20216 8676 20220 8732
rect 20156 8672 20220 8676
rect 20236 8732 20300 8736
rect 20236 8676 20240 8732
rect 20240 8676 20296 8732
rect 20296 8676 20300 8732
rect 20236 8672 20300 8676
rect 29518 8732 29582 8736
rect 29518 8676 29522 8732
rect 29522 8676 29578 8732
rect 29578 8676 29582 8732
rect 29518 8672 29582 8676
rect 29598 8732 29662 8736
rect 29598 8676 29602 8732
rect 29602 8676 29658 8732
rect 29658 8676 29662 8732
rect 29598 8672 29662 8676
rect 29678 8732 29742 8736
rect 29678 8676 29682 8732
rect 29682 8676 29738 8732
rect 29738 8676 29742 8732
rect 29678 8672 29742 8676
rect 29758 8732 29822 8736
rect 29758 8676 29762 8732
rect 29762 8676 29818 8732
rect 29818 8676 29822 8732
rect 29758 8672 29822 8676
rect 39040 8732 39104 8736
rect 39040 8676 39044 8732
rect 39044 8676 39100 8732
rect 39100 8676 39104 8732
rect 39040 8672 39104 8676
rect 39120 8732 39184 8736
rect 39120 8676 39124 8732
rect 39124 8676 39180 8732
rect 39180 8676 39184 8732
rect 39120 8672 39184 8676
rect 39200 8732 39264 8736
rect 39200 8676 39204 8732
rect 39204 8676 39260 8732
rect 39260 8676 39264 8732
rect 39200 8672 39264 8676
rect 39280 8732 39344 8736
rect 39280 8676 39284 8732
rect 39284 8676 39340 8732
rect 39340 8676 39344 8732
rect 39280 8672 39344 8676
rect 7052 8664 7116 8668
rect 7052 8608 7066 8664
rect 7066 8608 7116 8664
rect 7052 8604 7116 8608
rect 26188 8468 26252 8532
rect 28396 8604 28460 8668
rect 28580 8604 28644 8668
rect 5713 8188 5777 8192
rect 5713 8132 5717 8188
rect 5717 8132 5773 8188
rect 5773 8132 5777 8188
rect 5713 8128 5777 8132
rect 5793 8188 5857 8192
rect 5793 8132 5797 8188
rect 5797 8132 5853 8188
rect 5853 8132 5857 8188
rect 5793 8128 5857 8132
rect 5873 8188 5937 8192
rect 5873 8132 5877 8188
rect 5877 8132 5933 8188
rect 5933 8132 5937 8188
rect 5873 8128 5937 8132
rect 5953 8188 6017 8192
rect 5953 8132 5957 8188
rect 5957 8132 6013 8188
rect 6013 8132 6017 8188
rect 5953 8128 6017 8132
rect 3188 7924 3252 7988
rect 9444 8196 9508 8260
rect 15235 8188 15299 8192
rect 15235 8132 15239 8188
rect 15239 8132 15295 8188
rect 15295 8132 15299 8188
rect 15235 8128 15299 8132
rect 15315 8188 15379 8192
rect 15315 8132 15319 8188
rect 15319 8132 15375 8188
rect 15375 8132 15379 8188
rect 15315 8128 15379 8132
rect 15395 8188 15459 8192
rect 15395 8132 15399 8188
rect 15399 8132 15455 8188
rect 15455 8132 15459 8188
rect 15395 8128 15459 8132
rect 15475 8188 15539 8192
rect 15475 8132 15479 8188
rect 15479 8132 15535 8188
rect 15535 8132 15539 8188
rect 15475 8128 15539 8132
rect 13492 8060 13556 8124
rect 24757 8188 24821 8192
rect 24757 8132 24761 8188
rect 24761 8132 24817 8188
rect 24817 8132 24821 8188
rect 24757 8128 24821 8132
rect 24837 8188 24901 8192
rect 24837 8132 24841 8188
rect 24841 8132 24897 8188
rect 24897 8132 24901 8188
rect 24837 8128 24901 8132
rect 24917 8188 24981 8192
rect 24917 8132 24921 8188
rect 24921 8132 24977 8188
rect 24977 8132 24981 8188
rect 24917 8128 24981 8132
rect 24997 8188 25061 8192
rect 24997 8132 25001 8188
rect 25001 8132 25057 8188
rect 25057 8132 25061 8188
rect 24997 8128 25061 8132
rect 34279 8188 34343 8192
rect 34279 8132 34283 8188
rect 34283 8132 34339 8188
rect 34339 8132 34343 8188
rect 34279 8128 34343 8132
rect 34359 8188 34423 8192
rect 34359 8132 34363 8188
rect 34363 8132 34419 8188
rect 34419 8132 34423 8188
rect 34359 8128 34423 8132
rect 34439 8188 34503 8192
rect 34439 8132 34443 8188
rect 34443 8132 34499 8188
rect 34499 8132 34503 8188
rect 34439 8128 34503 8132
rect 34519 8188 34583 8192
rect 34519 8132 34523 8188
rect 34523 8132 34579 8188
rect 34579 8132 34583 8188
rect 34519 8128 34583 8132
rect 29132 8060 29196 8124
rect 24532 7924 24596 7988
rect 23428 7652 23492 7716
rect 10474 7644 10538 7648
rect 10474 7588 10478 7644
rect 10478 7588 10534 7644
rect 10534 7588 10538 7644
rect 10474 7584 10538 7588
rect 10554 7644 10618 7648
rect 10554 7588 10558 7644
rect 10558 7588 10614 7644
rect 10614 7588 10618 7644
rect 10554 7584 10618 7588
rect 10634 7644 10698 7648
rect 10634 7588 10638 7644
rect 10638 7588 10694 7644
rect 10694 7588 10698 7644
rect 10634 7584 10698 7588
rect 10714 7644 10778 7648
rect 10714 7588 10718 7644
rect 10718 7588 10774 7644
rect 10774 7588 10778 7644
rect 10714 7584 10778 7588
rect 19996 7644 20060 7648
rect 19996 7588 20000 7644
rect 20000 7588 20056 7644
rect 20056 7588 20060 7644
rect 19996 7584 20060 7588
rect 20076 7644 20140 7648
rect 20076 7588 20080 7644
rect 20080 7588 20136 7644
rect 20136 7588 20140 7644
rect 20076 7584 20140 7588
rect 20156 7644 20220 7648
rect 20156 7588 20160 7644
rect 20160 7588 20216 7644
rect 20216 7588 20220 7644
rect 20156 7584 20220 7588
rect 20236 7644 20300 7648
rect 20236 7588 20240 7644
rect 20240 7588 20296 7644
rect 20296 7588 20300 7644
rect 20236 7584 20300 7588
rect 29518 7644 29582 7648
rect 29518 7588 29522 7644
rect 29522 7588 29578 7644
rect 29578 7588 29582 7644
rect 29518 7584 29582 7588
rect 29598 7644 29662 7648
rect 29598 7588 29602 7644
rect 29602 7588 29658 7644
rect 29658 7588 29662 7644
rect 29598 7584 29662 7588
rect 29678 7644 29742 7648
rect 29678 7588 29682 7644
rect 29682 7588 29738 7644
rect 29738 7588 29742 7644
rect 29678 7584 29742 7588
rect 29758 7644 29822 7648
rect 29758 7588 29762 7644
rect 29762 7588 29818 7644
rect 29818 7588 29822 7644
rect 29758 7584 29822 7588
rect 39040 7644 39104 7648
rect 39040 7588 39044 7644
rect 39044 7588 39100 7644
rect 39100 7588 39104 7644
rect 39040 7584 39104 7588
rect 39120 7644 39184 7648
rect 39120 7588 39124 7644
rect 39124 7588 39180 7644
rect 39180 7588 39184 7644
rect 39120 7584 39184 7588
rect 39200 7644 39264 7648
rect 39200 7588 39204 7644
rect 39204 7588 39260 7644
rect 39260 7588 39264 7644
rect 39200 7584 39264 7588
rect 39280 7644 39344 7648
rect 39280 7588 39284 7644
rect 39284 7588 39340 7644
rect 39340 7588 39344 7644
rect 39280 7584 39344 7588
rect 5713 7100 5777 7104
rect 5713 7044 5717 7100
rect 5717 7044 5773 7100
rect 5773 7044 5777 7100
rect 5713 7040 5777 7044
rect 5793 7100 5857 7104
rect 5793 7044 5797 7100
rect 5797 7044 5853 7100
rect 5853 7044 5857 7100
rect 5793 7040 5857 7044
rect 5873 7100 5937 7104
rect 5873 7044 5877 7100
rect 5877 7044 5933 7100
rect 5933 7044 5937 7100
rect 5873 7040 5937 7044
rect 5953 7100 6017 7104
rect 5953 7044 5957 7100
rect 5957 7044 6013 7100
rect 6013 7044 6017 7100
rect 5953 7040 6017 7044
rect 15235 7100 15299 7104
rect 15235 7044 15239 7100
rect 15239 7044 15295 7100
rect 15295 7044 15299 7100
rect 15235 7040 15299 7044
rect 15315 7100 15379 7104
rect 15315 7044 15319 7100
rect 15319 7044 15375 7100
rect 15375 7044 15379 7100
rect 15315 7040 15379 7044
rect 15395 7100 15459 7104
rect 15395 7044 15399 7100
rect 15399 7044 15455 7100
rect 15455 7044 15459 7100
rect 15395 7040 15459 7044
rect 15475 7100 15539 7104
rect 15475 7044 15479 7100
rect 15479 7044 15535 7100
rect 15535 7044 15539 7100
rect 15475 7040 15539 7044
rect 24757 7100 24821 7104
rect 24757 7044 24761 7100
rect 24761 7044 24817 7100
rect 24817 7044 24821 7100
rect 24757 7040 24821 7044
rect 24837 7100 24901 7104
rect 24837 7044 24841 7100
rect 24841 7044 24897 7100
rect 24897 7044 24901 7100
rect 24837 7040 24901 7044
rect 24917 7100 24981 7104
rect 24917 7044 24921 7100
rect 24921 7044 24977 7100
rect 24977 7044 24981 7100
rect 24917 7040 24981 7044
rect 24997 7100 25061 7104
rect 24997 7044 25001 7100
rect 25001 7044 25057 7100
rect 25057 7044 25061 7100
rect 24997 7040 25061 7044
rect 34279 7100 34343 7104
rect 34279 7044 34283 7100
rect 34283 7044 34339 7100
rect 34339 7044 34343 7100
rect 34279 7040 34343 7044
rect 34359 7100 34423 7104
rect 34359 7044 34363 7100
rect 34363 7044 34419 7100
rect 34419 7044 34423 7100
rect 34359 7040 34423 7044
rect 34439 7100 34503 7104
rect 34439 7044 34443 7100
rect 34443 7044 34499 7100
rect 34499 7044 34503 7100
rect 34439 7040 34503 7044
rect 34519 7100 34583 7104
rect 34519 7044 34523 7100
rect 34523 7044 34579 7100
rect 34579 7044 34583 7100
rect 34519 7040 34583 7044
rect 12572 6972 12636 7036
rect 4108 6836 4172 6900
rect 31156 6836 31220 6900
rect 6500 6760 6564 6764
rect 6500 6704 6514 6760
rect 6514 6704 6564 6760
rect 6500 6700 6564 6704
rect 7052 6700 7116 6764
rect 9628 6700 9692 6764
rect 15700 6700 15764 6764
rect 22324 6624 22388 6628
rect 22324 6568 22374 6624
rect 22374 6568 22388 6624
rect 22324 6564 22388 6568
rect 10474 6556 10538 6560
rect 10474 6500 10478 6556
rect 10478 6500 10534 6556
rect 10534 6500 10538 6556
rect 10474 6496 10538 6500
rect 10554 6556 10618 6560
rect 10554 6500 10558 6556
rect 10558 6500 10614 6556
rect 10614 6500 10618 6556
rect 10554 6496 10618 6500
rect 10634 6556 10698 6560
rect 10634 6500 10638 6556
rect 10638 6500 10694 6556
rect 10694 6500 10698 6556
rect 10634 6496 10698 6500
rect 10714 6556 10778 6560
rect 10714 6500 10718 6556
rect 10718 6500 10774 6556
rect 10774 6500 10778 6556
rect 10714 6496 10778 6500
rect 19996 6556 20060 6560
rect 19996 6500 20000 6556
rect 20000 6500 20056 6556
rect 20056 6500 20060 6556
rect 19996 6496 20060 6500
rect 20076 6556 20140 6560
rect 20076 6500 20080 6556
rect 20080 6500 20136 6556
rect 20136 6500 20140 6556
rect 20076 6496 20140 6500
rect 20156 6556 20220 6560
rect 20156 6500 20160 6556
rect 20160 6500 20216 6556
rect 20216 6500 20220 6556
rect 20156 6496 20220 6500
rect 20236 6556 20300 6560
rect 20236 6500 20240 6556
rect 20240 6500 20296 6556
rect 20296 6500 20300 6556
rect 20236 6496 20300 6500
rect 29518 6556 29582 6560
rect 29518 6500 29522 6556
rect 29522 6500 29578 6556
rect 29578 6500 29582 6556
rect 29518 6496 29582 6500
rect 29598 6556 29662 6560
rect 29598 6500 29602 6556
rect 29602 6500 29658 6556
rect 29658 6500 29662 6556
rect 29598 6496 29662 6500
rect 29678 6556 29742 6560
rect 29678 6500 29682 6556
rect 29682 6500 29738 6556
rect 29738 6500 29742 6556
rect 29678 6496 29742 6500
rect 29758 6556 29822 6560
rect 29758 6500 29762 6556
rect 29762 6500 29818 6556
rect 29818 6500 29822 6556
rect 29758 6496 29822 6500
rect 39040 6556 39104 6560
rect 39040 6500 39044 6556
rect 39044 6500 39100 6556
rect 39100 6500 39104 6556
rect 39040 6496 39104 6500
rect 39120 6556 39184 6560
rect 39120 6500 39124 6556
rect 39124 6500 39180 6556
rect 39180 6500 39184 6556
rect 39120 6496 39184 6500
rect 39200 6556 39264 6560
rect 39200 6500 39204 6556
rect 39204 6500 39260 6556
rect 39260 6500 39264 6556
rect 39200 6496 39264 6500
rect 39280 6556 39344 6560
rect 39280 6500 39284 6556
rect 39284 6500 39340 6556
rect 39340 6500 39344 6556
rect 39280 6496 39344 6500
rect 13860 6428 13924 6492
rect 26924 6428 26988 6492
rect 19564 6292 19628 6356
rect 25820 6292 25884 6356
rect 5713 6012 5777 6016
rect 5713 5956 5717 6012
rect 5717 5956 5773 6012
rect 5773 5956 5777 6012
rect 5713 5952 5777 5956
rect 5793 6012 5857 6016
rect 5793 5956 5797 6012
rect 5797 5956 5853 6012
rect 5853 5956 5857 6012
rect 5793 5952 5857 5956
rect 5873 6012 5937 6016
rect 5873 5956 5877 6012
rect 5877 5956 5933 6012
rect 5933 5956 5937 6012
rect 5873 5952 5937 5956
rect 5953 6012 6017 6016
rect 5953 5956 5957 6012
rect 5957 5956 6013 6012
rect 6013 5956 6017 6012
rect 5953 5952 6017 5956
rect 25820 6020 25884 6084
rect 15235 6012 15299 6016
rect 15235 5956 15239 6012
rect 15239 5956 15295 6012
rect 15295 5956 15299 6012
rect 15235 5952 15299 5956
rect 15315 6012 15379 6016
rect 15315 5956 15319 6012
rect 15319 5956 15375 6012
rect 15375 5956 15379 6012
rect 15315 5952 15379 5956
rect 15395 6012 15459 6016
rect 15395 5956 15399 6012
rect 15399 5956 15455 6012
rect 15455 5956 15459 6012
rect 15395 5952 15459 5956
rect 15475 6012 15539 6016
rect 15475 5956 15479 6012
rect 15479 5956 15535 6012
rect 15535 5956 15539 6012
rect 15475 5952 15539 5956
rect 24757 6012 24821 6016
rect 24757 5956 24761 6012
rect 24761 5956 24817 6012
rect 24817 5956 24821 6012
rect 24757 5952 24821 5956
rect 24837 6012 24901 6016
rect 24837 5956 24841 6012
rect 24841 5956 24897 6012
rect 24897 5956 24901 6012
rect 24837 5952 24901 5956
rect 24917 6012 24981 6016
rect 24917 5956 24921 6012
rect 24921 5956 24977 6012
rect 24977 5956 24981 6012
rect 24917 5952 24981 5956
rect 24997 6012 25061 6016
rect 24997 5956 25001 6012
rect 25001 5956 25057 6012
rect 25057 5956 25061 6012
rect 24997 5952 25061 5956
rect 34279 6012 34343 6016
rect 34279 5956 34283 6012
rect 34283 5956 34339 6012
rect 34339 5956 34343 6012
rect 34279 5952 34343 5956
rect 34359 6012 34423 6016
rect 34359 5956 34363 6012
rect 34363 5956 34419 6012
rect 34419 5956 34423 6012
rect 34359 5952 34423 5956
rect 34439 6012 34503 6016
rect 34439 5956 34443 6012
rect 34443 5956 34499 6012
rect 34499 5956 34503 6012
rect 34439 5952 34503 5956
rect 34519 6012 34583 6016
rect 34519 5956 34523 6012
rect 34523 5956 34579 6012
rect 34579 5956 34583 6012
rect 34519 5952 34583 5956
rect 25636 5944 25700 5948
rect 25636 5888 25650 5944
rect 25650 5888 25700 5944
rect 25636 5884 25700 5888
rect 26188 5884 26252 5948
rect 30420 5884 30484 5948
rect 8892 5612 8956 5676
rect 9628 5672 9692 5676
rect 9628 5616 9678 5672
rect 9678 5616 9692 5672
rect 9628 5612 9692 5616
rect 11100 5612 11164 5676
rect 15884 5476 15948 5540
rect 16620 5536 16684 5540
rect 16620 5480 16670 5536
rect 16670 5480 16684 5536
rect 16620 5476 16684 5480
rect 10474 5468 10538 5472
rect 10474 5412 10478 5468
rect 10478 5412 10534 5468
rect 10534 5412 10538 5468
rect 10474 5408 10538 5412
rect 10554 5468 10618 5472
rect 10554 5412 10558 5468
rect 10558 5412 10614 5468
rect 10614 5412 10618 5468
rect 10554 5408 10618 5412
rect 10634 5468 10698 5472
rect 10634 5412 10638 5468
rect 10638 5412 10694 5468
rect 10694 5412 10698 5468
rect 10634 5408 10698 5412
rect 10714 5468 10778 5472
rect 10714 5412 10718 5468
rect 10718 5412 10774 5468
rect 10774 5412 10778 5468
rect 10714 5408 10778 5412
rect 19996 5468 20060 5472
rect 19996 5412 20000 5468
rect 20000 5412 20056 5468
rect 20056 5412 20060 5468
rect 19996 5408 20060 5412
rect 20076 5468 20140 5472
rect 20076 5412 20080 5468
rect 20080 5412 20136 5468
rect 20136 5412 20140 5468
rect 20076 5408 20140 5412
rect 20156 5468 20220 5472
rect 20156 5412 20160 5468
rect 20160 5412 20216 5468
rect 20216 5412 20220 5468
rect 20156 5408 20220 5412
rect 20236 5468 20300 5472
rect 20236 5412 20240 5468
rect 20240 5412 20296 5468
rect 20296 5412 20300 5468
rect 20236 5408 20300 5412
rect 6316 5340 6380 5404
rect 13308 5340 13372 5404
rect 2820 5204 2884 5268
rect 28212 5204 28276 5268
rect 33732 5476 33796 5540
rect 29518 5468 29582 5472
rect 29518 5412 29522 5468
rect 29522 5412 29578 5468
rect 29578 5412 29582 5468
rect 29518 5408 29582 5412
rect 29598 5468 29662 5472
rect 29598 5412 29602 5468
rect 29602 5412 29658 5468
rect 29658 5412 29662 5468
rect 29598 5408 29662 5412
rect 29678 5468 29742 5472
rect 29678 5412 29682 5468
rect 29682 5412 29738 5468
rect 29738 5412 29742 5468
rect 29678 5408 29742 5412
rect 29758 5468 29822 5472
rect 29758 5412 29762 5468
rect 29762 5412 29818 5468
rect 29818 5412 29822 5468
rect 29758 5408 29822 5412
rect 39040 5468 39104 5472
rect 39040 5412 39044 5468
rect 39044 5412 39100 5468
rect 39100 5412 39104 5468
rect 39040 5408 39104 5412
rect 39120 5468 39184 5472
rect 39120 5412 39124 5468
rect 39124 5412 39180 5468
rect 39180 5412 39184 5468
rect 39120 5408 39184 5412
rect 39200 5468 39264 5472
rect 39200 5412 39204 5468
rect 39204 5412 39260 5468
rect 39260 5412 39264 5468
rect 39200 5408 39264 5412
rect 39280 5468 39344 5472
rect 39280 5412 39284 5468
rect 39284 5412 39340 5468
rect 39340 5412 39344 5468
rect 39280 5408 39344 5412
rect 7604 4932 7668 4996
rect 5713 4924 5777 4928
rect 5713 4868 5717 4924
rect 5717 4868 5773 4924
rect 5773 4868 5777 4924
rect 5713 4864 5777 4868
rect 5793 4924 5857 4928
rect 5793 4868 5797 4924
rect 5797 4868 5853 4924
rect 5853 4868 5857 4924
rect 5793 4864 5857 4868
rect 5873 4924 5937 4928
rect 5873 4868 5877 4924
rect 5877 4868 5933 4924
rect 5933 4868 5937 4924
rect 5873 4864 5937 4868
rect 5953 4924 6017 4928
rect 5953 4868 5957 4924
rect 5957 4868 6013 4924
rect 6013 4868 6017 4924
rect 5953 4864 6017 4868
rect 15235 4924 15299 4928
rect 15235 4868 15239 4924
rect 15239 4868 15295 4924
rect 15295 4868 15299 4924
rect 15235 4864 15299 4868
rect 15315 4924 15379 4928
rect 15315 4868 15319 4924
rect 15319 4868 15375 4924
rect 15375 4868 15379 4924
rect 15315 4864 15379 4868
rect 15395 4924 15459 4928
rect 15395 4868 15399 4924
rect 15399 4868 15455 4924
rect 15455 4868 15459 4924
rect 15395 4864 15459 4868
rect 15475 4924 15539 4928
rect 15475 4868 15479 4924
rect 15479 4868 15535 4924
rect 15535 4868 15539 4924
rect 15475 4864 15539 4868
rect 24757 4924 24821 4928
rect 24757 4868 24761 4924
rect 24761 4868 24817 4924
rect 24817 4868 24821 4924
rect 24757 4864 24821 4868
rect 24837 4924 24901 4928
rect 24837 4868 24841 4924
rect 24841 4868 24897 4924
rect 24897 4868 24901 4924
rect 24837 4864 24901 4868
rect 24917 4924 24981 4928
rect 24917 4868 24921 4924
rect 24921 4868 24977 4924
rect 24977 4868 24981 4924
rect 24917 4864 24981 4868
rect 24997 4924 25061 4928
rect 24997 4868 25001 4924
rect 25001 4868 25057 4924
rect 25057 4868 25061 4924
rect 24997 4864 25061 4868
rect 34279 4924 34343 4928
rect 34279 4868 34283 4924
rect 34283 4868 34339 4924
rect 34339 4868 34343 4924
rect 34279 4864 34343 4868
rect 34359 4924 34423 4928
rect 34359 4868 34363 4924
rect 34363 4868 34419 4924
rect 34419 4868 34423 4924
rect 34359 4864 34423 4868
rect 34439 4924 34503 4928
rect 34439 4868 34443 4924
rect 34443 4868 34499 4924
rect 34499 4868 34503 4924
rect 34439 4864 34503 4868
rect 34519 4924 34583 4928
rect 34519 4868 34523 4924
rect 34523 4868 34579 4924
rect 34579 4868 34583 4924
rect 34519 4864 34583 4868
rect 13308 4856 13372 4860
rect 13308 4800 13358 4856
rect 13358 4800 13372 4856
rect 13308 4796 13372 4800
rect 27108 4388 27172 4452
rect 10474 4380 10538 4384
rect 10474 4324 10478 4380
rect 10478 4324 10534 4380
rect 10534 4324 10538 4380
rect 10474 4320 10538 4324
rect 10554 4380 10618 4384
rect 10554 4324 10558 4380
rect 10558 4324 10614 4380
rect 10614 4324 10618 4380
rect 10554 4320 10618 4324
rect 10634 4380 10698 4384
rect 10634 4324 10638 4380
rect 10638 4324 10694 4380
rect 10694 4324 10698 4380
rect 10634 4320 10698 4324
rect 10714 4380 10778 4384
rect 10714 4324 10718 4380
rect 10718 4324 10774 4380
rect 10774 4324 10778 4380
rect 10714 4320 10778 4324
rect 19996 4380 20060 4384
rect 19996 4324 20000 4380
rect 20000 4324 20056 4380
rect 20056 4324 20060 4380
rect 19996 4320 20060 4324
rect 20076 4380 20140 4384
rect 20076 4324 20080 4380
rect 20080 4324 20136 4380
rect 20136 4324 20140 4380
rect 20076 4320 20140 4324
rect 20156 4380 20220 4384
rect 20156 4324 20160 4380
rect 20160 4324 20216 4380
rect 20216 4324 20220 4380
rect 20156 4320 20220 4324
rect 20236 4380 20300 4384
rect 20236 4324 20240 4380
rect 20240 4324 20296 4380
rect 20296 4324 20300 4380
rect 20236 4320 20300 4324
rect 5212 4116 5276 4180
rect 29518 4380 29582 4384
rect 29518 4324 29522 4380
rect 29522 4324 29578 4380
rect 29578 4324 29582 4380
rect 29518 4320 29582 4324
rect 29598 4380 29662 4384
rect 29598 4324 29602 4380
rect 29602 4324 29658 4380
rect 29658 4324 29662 4380
rect 29598 4320 29662 4324
rect 29678 4380 29742 4384
rect 29678 4324 29682 4380
rect 29682 4324 29738 4380
rect 29738 4324 29742 4380
rect 29678 4320 29742 4324
rect 29758 4380 29822 4384
rect 29758 4324 29762 4380
rect 29762 4324 29818 4380
rect 29818 4324 29822 4380
rect 29758 4320 29822 4324
rect 39040 4380 39104 4384
rect 39040 4324 39044 4380
rect 39044 4324 39100 4380
rect 39100 4324 39104 4380
rect 39040 4320 39104 4324
rect 39120 4380 39184 4384
rect 39120 4324 39124 4380
rect 39124 4324 39180 4380
rect 39180 4324 39184 4380
rect 39120 4320 39184 4324
rect 39200 4380 39264 4384
rect 39200 4324 39204 4380
rect 39204 4324 39260 4380
rect 39260 4324 39264 4380
rect 39200 4320 39264 4324
rect 39280 4380 39344 4384
rect 39280 4324 39284 4380
rect 39284 4324 39340 4380
rect 39340 4324 39344 4380
rect 39280 4320 39344 4324
rect 12204 4040 12268 4044
rect 12204 3984 12254 4040
rect 12254 3984 12268 4040
rect 5713 3836 5777 3840
rect 5713 3780 5717 3836
rect 5717 3780 5773 3836
rect 5773 3780 5777 3836
rect 5713 3776 5777 3780
rect 5793 3836 5857 3840
rect 5793 3780 5797 3836
rect 5797 3780 5853 3836
rect 5853 3780 5857 3836
rect 5793 3776 5857 3780
rect 5873 3836 5937 3840
rect 5873 3780 5877 3836
rect 5877 3780 5933 3836
rect 5933 3780 5937 3836
rect 5873 3776 5937 3780
rect 5953 3836 6017 3840
rect 5953 3780 5957 3836
rect 5957 3780 6013 3836
rect 6013 3780 6017 3836
rect 5953 3776 6017 3780
rect 3188 3572 3252 3636
rect 12204 3980 12268 3984
rect 17908 4040 17972 4044
rect 17908 3984 17958 4040
rect 17958 3984 17972 4040
rect 12020 3844 12084 3908
rect 17908 3980 17972 3984
rect 18276 4040 18340 4044
rect 18276 3984 18290 4040
rect 18290 3984 18340 4040
rect 18276 3980 18340 3984
rect 30052 4040 30116 4044
rect 30052 3984 30066 4040
rect 30066 3984 30116 4040
rect 30052 3980 30116 3984
rect 32628 3904 32692 3908
rect 32628 3848 32678 3904
rect 32678 3848 32692 3904
rect 32628 3844 32692 3848
rect 15235 3836 15299 3840
rect 15235 3780 15239 3836
rect 15239 3780 15295 3836
rect 15295 3780 15299 3836
rect 15235 3776 15299 3780
rect 15315 3836 15379 3840
rect 15315 3780 15319 3836
rect 15319 3780 15375 3836
rect 15375 3780 15379 3836
rect 15315 3776 15379 3780
rect 15395 3836 15459 3840
rect 15395 3780 15399 3836
rect 15399 3780 15455 3836
rect 15455 3780 15459 3836
rect 15395 3776 15459 3780
rect 15475 3836 15539 3840
rect 15475 3780 15479 3836
rect 15479 3780 15535 3836
rect 15535 3780 15539 3836
rect 15475 3776 15539 3780
rect 24757 3836 24821 3840
rect 24757 3780 24761 3836
rect 24761 3780 24817 3836
rect 24817 3780 24821 3836
rect 24757 3776 24821 3780
rect 24837 3836 24901 3840
rect 24837 3780 24841 3836
rect 24841 3780 24897 3836
rect 24897 3780 24901 3836
rect 24837 3776 24901 3780
rect 24917 3836 24981 3840
rect 24917 3780 24921 3836
rect 24921 3780 24977 3836
rect 24977 3780 24981 3836
rect 24917 3776 24981 3780
rect 24997 3836 25061 3840
rect 24997 3780 25001 3836
rect 25001 3780 25057 3836
rect 25057 3780 25061 3836
rect 24997 3776 25061 3780
rect 34279 3836 34343 3840
rect 34279 3780 34283 3836
rect 34283 3780 34339 3836
rect 34339 3780 34343 3836
rect 34279 3776 34343 3780
rect 34359 3836 34423 3840
rect 34359 3780 34363 3836
rect 34363 3780 34419 3836
rect 34419 3780 34423 3836
rect 34359 3776 34423 3780
rect 34439 3836 34503 3840
rect 34439 3780 34443 3836
rect 34443 3780 34499 3836
rect 34499 3780 34503 3836
rect 34439 3776 34503 3780
rect 34519 3836 34583 3840
rect 34519 3780 34523 3836
rect 34523 3780 34579 3836
rect 34579 3780 34583 3836
rect 34519 3776 34583 3780
rect 28948 3300 29012 3364
rect 34652 3300 34716 3364
rect 10474 3292 10538 3296
rect 10474 3236 10478 3292
rect 10478 3236 10534 3292
rect 10534 3236 10538 3292
rect 10474 3232 10538 3236
rect 10554 3292 10618 3296
rect 10554 3236 10558 3292
rect 10558 3236 10614 3292
rect 10614 3236 10618 3292
rect 10554 3232 10618 3236
rect 10634 3292 10698 3296
rect 10634 3236 10638 3292
rect 10638 3236 10694 3292
rect 10694 3236 10698 3292
rect 10634 3232 10698 3236
rect 10714 3292 10778 3296
rect 10714 3236 10718 3292
rect 10718 3236 10774 3292
rect 10774 3236 10778 3292
rect 10714 3232 10778 3236
rect 19996 3292 20060 3296
rect 19996 3236 20000 3292
rect 20000 3236 20056 3292
rect 20056 3236 20060 3292
rect 19996 3232 20060 3236
rect 20076 3292 20140 3296
rect 20076 3236 20080 3292
rect 20080 3236 20136 3292
rect 20136 3236 20140 3292
rect 20076 3232 20140 3236
rect 20156 3292 20220 3296
rect 20156 3236 20160 3292
rect 20160 3236 20216 3292
rect 20216 3236 20220 3292
rect 20156 3232 20220 3236
rect 20236 3292 20300 3296
rect 20236 3236 20240 3292
rect 20240 3236 20296 3292
rect 20296 3236 20300 3292
rect 20236 3232 20300 3236
rect 29518 3292 29582 3296
rect 29518 3236 29522 3292
rect 29522 3236 29578 3292
rect 29578 3236 29582 3292
rect 29518 3232 29582 3236
rect 29598 3292 29662 3296
rect 29598 3236 29602 3292
rect 29602 3236 29658 3292
rect 29658 3236 29662 3292
rect 29598 3232 29662 3236
rect 29678 3292 29742 3296
rect 29678 3236 29682 3292
rect 29682 3236 29738 3292
rect 29738 3236 29742 3292
rect 29678 3232 29742 3236
rect 29758 3292 29822 3296
rect 29758 3236 29762 3292
rect 29762 3236 29818 3292
rect 29818 3236 29822 3292
rect 29758 3232 29822 3236
rect 39040 3292 39104 3296
rect 39040 3236 39044 3292
rect 39044 3236 39100 3292
rect 39100 3236 39104 3292
rect 39040 3232 39104 3236
rect 39120 3292 39184 3296
rect 39120 3236 39124 3292
rect 39124 3236 39180 3292
rect 39180 3236 39184 3292
rect 39120 3232 39184 3236
rect 39200 3292 39264 3296
rect 39200 3236 39204 3292
rect 39204 3236 39260 3292
rect 39260 3236 39264 3292
rect 39200 3232 39264 3236
rect 39280 3292 39344 3296
rect 39280 3236 39284 3292
rect 39284 3236 39340 3292
rect 39340 3236 39344 3292
rect 39280 3232 39344 3236
rect 14044 3088 14108 3092
rect 14044 3032 14094 3088
rect 14094 3032 14108 3088
rect 14044 3028 14108 3032
rect 26740 3164 26804 3228
rect 5713 2748 5777 2752
rect 5713 2692 5717 2748
rect 5717 2692 5773 2748
rect 5773 2692 5777 2748
rect 5713 2688 5777 2692
rect 5793 2748 5857 2752
rect 5793 2692 5797 2748
rect 5797 2692 5853 2748
rect 5853 2692 5857 2748
rect 5793 2688 5857 2692
rect 5873 2748 5937 2752
rect 5873 2692 5877 2748
rect 5877 2692 5933 2748
rect 5933 2692 5937 2748
rect 5873 2688 5937 2692
rect 5953 2748 6017 2752
rect 5953 2692 5957 2748
rect 5957 2692 6013 2748
rect 6013 2692 6017 2748
rect 5953 2688 6017 2692
rect 15235 2748 15299 2752
rect 15235 2692 15239 2748
rect 15239 2692 15295 2748
rect 15295 2692 15299 2748
rect 15235 2688 15299 2692
rect 15315 2748 15379 2752
rect 15315 2692 15319 2748
rect 15319 2692 15375 2748
rect 15375 2692 15379 2748
rect 15315 2688 15379 2692
rect 15395 2748 15459 2752
rect 15395 2692 15399 2748
rect 15399 2692 15455 2748
rect 15455 2692 15459 2748
rect 15395 2688 15459 2692
rect 15475 2748 15539 2752
rect 15475 2692 15479 2748
rect 15479 2692 15535 2748
rect 15535 2692 15539 2748
rect 15475 2688 15539 2692
rect 24757 2748 24821 2752
rect 24757 2692 24761 2748
rect 24761 2692 24817 2748
rect 24817 2692 24821 2748
rect 24757 2688 24821 2692
rect 24837 2748 24901 2752
rect 24837 2692 24841 2748
rect 24841 2692 24897 2748
rect 24897 2692 24901 2748
rect 24837 2688 24901 2692
rect 24917 2748 24981 2752
rect 24917 2692 24921 2748
rect 24921 2692 24977 2748
rect 24977 2692 24981 2748
rect 24917 2688 24981 2692
rect 24997 2748 25061 2752
rect 24997 2692 25001 2748
rect 25001 2692 25057 2748
rect 25057 2692 25061 2748
rect 24997 2688 25061 2692
rect 34279 2748 34343 2752
rect 34279 2692 34283 2748
rect 34283 2692 34339 2748
rect 34339 2692 34343 2748
rect 34279 2688 34343 2692
rect 34359 2748 34423 2752
rect 34359 2692 34363 2748
rect 34363 2692 34419 2748
rect 34419 2692 34423 2748
rect 34359 2688 34423 2692
rect 34439 2748 34503 2752
rect 34439 2692 34443 2748
rect 34443 2692 34499 2748
rect 34499 2692 34503 2748
rect 34439 2688 34503 2692
rect 34519 2748 34583 2752
rect 34519 2692 34523 2748
rect 34523 2692 34579 2748
rect 34579 2692 34583 2748
rect 34519 2688 34583 2692
rect 17172 2680 17236 2684
rect 17172 2624 17186 2680
rect 17186 2624 17236 2680
rect 17172 2620 17236 2624
rect 27660 2620 27724 2684
rect 33180 2680 33244 2684
rect 33180 2624 33230 2680
rect 33230 2624 33244 2680
rect 33180 2620 33244 2624
rect 5396 2484 5460 2548
rect 23980 2484 24044 2548
rect 10474 2204 10538 2208
rect 10474 2148 10478 2204
rect 10478 2148 10534 2204
rect 10534 2148 10538 2204
rect 10474 2144 10538 2148
rect 10554 2204 10618 2208
rect 10554 2148 10558 2204
rect 10558 2148 10614 2204
rect 10614 2148 10618 2204
rect 10554 2144 10618 2148
rect 10634 2204 10698 2208
rect 10634 2148 10638 2204
rect 10638 2148 10694 2204
rect 10694 2148 10698 2204
rect 10634 2144 10698 2148
rect 10714 2204 10778 2208
rect 10714 2148 10718 2204
rect 10718 2148 10774 2204
rect 10774 2148 10778 2204
rect 10714 2144 10778 2148
rect 19996 2204 20060 2208
rect 19996 2148 20000 2204
rect 20000 2148 20056 2204
rect 20056 2148 20060 2204
rect 19996 2144 20060 2148
rect 20076 2204 20140 2208
rect 20076 2148 20080 2204
rect 20080 2148 20136 2204
rect 20136 2148 20140 2204
rect 20076 2144 20140 2148
rect 20156 2204 20220 2208
rect 20156 2148 20160 2204
rect 20160 2148 20216 2204
rect 20216 2148 20220 2204
rect 20156 2144 20220 2148
rect 20236 2204 20300 2208
rect 20236 2148 20240 2204
rect 20240 2148 20296 2204
rect 20296 2148 20300 2204
rect 20236 2144 20300 2148
rect 29518 2204 29582 2208
rect 29518 2148 29522 2204
rect 29522 2148 29578 2204
rect 29578 2148 29582 2204
rect 29518 2144 29582 2148
rect 29598 2204 29662 2208
rect 29598 2148 29602 2204
rect 29602 2148 29658 2204
rect 29658 2148 29662 2204
rect 29598 2144 29662 2148
rect 29678 2204 29742 2208
rect 29678 2148 29682 2204
rect 29682 2148 29738 2204
rect 29738 2148 29742 2204
rect 29678 2144 29742 2148
rect 29758 2204 29822 2208
rect 29758 2148 29762 2204
rect 29762 2148 29818 2204
rect 29818 2148 29822 2204
rect 29758 2144 29822 2148
rect 39040 2204 39104 2208
rect 39040 2148 39044 2204
rect 39044 2148 39100 2204
rect 39100 2148 39104 2204
rect 39040 2144 39104 2148
rect 39120 2204 39184 2208
rect 39120 2148 39124 2204
rect 39124 2148 39180 2204
rect 39180 2148 39184 2204
rect 39120 2144 39184 2148
rect 39200 2204 39264 2208
rect 39200 2148 39204 2204
rect 39204 2148 39260 2204
rect 39260 2148 39264 2204
rect 39200 2144 39264 2148
rect 39280 2204 39344 2208
rect 39280 2148 39284 2204
rect 39284 2148 39340 2204
rect 39340 2148 39344 2204
rect 39280 2144 39344 2148
rect 10180 1804 10244 1868
rect 2636 1260 2700 1324
<< metal4 >>
rect 5705 26688 6025 26704
rect 5705 26624 5713 26688
rect 5777 26624 5793 26688
rect 5857 26624 5873 26688
rect 5937 26624 5953 26688
rect 6017 26624 6025 26688
rect 5705 25600 6025 26624
rect 6315 26348 6381 26349
rect 6315 26284 6316 26348
rect 6380 26284 6381 26348
rect 6315 26283 6381 26284
rect 5705 25536 5713 25600
rect 5777 25536 5793 25600
rect 5857 25536 5873 25600
rect 5937 25536 5953 25600
rect 6017 25536 6025 25600
rect 5705 24512 6025 25536
rect 5705 24448 5713 24512
rect 5777 24448 5793 24512
rect 5857 24448 5873 24512
rect 5937 24448 5953 24512
rect 6017 24448 6025 24512
rect 5705 23424 6025 24448
rect 5705 23360 5713 23424
rect 5777 23360 5793 23424
rect 5857 23360 5873 23424
rect 5937 23360 5953 23424
rect 6017 23360 6025 23424
rect 5705 22336 6025 23360
rect 5705 22272 5713 22336
rect 5777 22272 5793 22336
rect 5857 22272 5873 22336
rect 5937 22272 5953 22336
rect 6017 22272 6025 22336
rect 5705 21248 6025 22272
rect 5705 21184 5713 21248
rect 5777 21184 5793 21248
rect 5857 21184 5873 21248
rect 5937 21184 5953 21248
rect 6017 21184 6025 21248
rect 5705 20160 6025 21184
rect 5705 20096 5713 20160
rect 5777 20096 5793 20160
rect 5857 20096 5873 20160
rect 5937 20096 5953 20160
rect 6017 20096 6025 20160
rect 5705 19072 6025 20096
rect 5705 19008 5713 19072
rect 5777 19008 5793 19072
rect 5857 19008 5873 19072
rect 5937 19008 5953 19072
rect 6017 19008 6025 19072
rect 5705 17984 6025 19008
rect 5705 17920 5713 17984
rect 5777 17920 5793 17984
rect 5857 17920 5873 17984
rect 5937 17920 5953 17984
rect 6017 17920 6025 17984
rect 5211 17100 5277 17101
rect 5211 17036 5212 17100
rect 5276 17036 5277 17100
rect 5211 17035 5277 17036
rect 2819 16692 2885 16693
rect 2819 16628 2820 16692
rect 2884 16628 2885 16692
rect 2819 16627 2885 16628
rect 2635 9756 2701 9757
rect 2635 9692 2636 9756
rect 2700 9692 2701 9756
rect 2635 9691 2701 9692
rect 2638 1325 2698 9691
rect 2822 5269 2882 16627
rect 3187 15332 3253 15333
rect 3187 15268 3188 15332
rect 3252 15268 3253 15332
rect 3187 15267 3253 15268
rect 4107 15332 4173 15333
rect 4107 15268 4108 15332
rect 4172 15268 4173 15332
rect 4107 15267 4173 15268
rect 3190 7989 3250 15267
rect 3187 7988 3253 7989
rect 3187 7924 3188 7988
rect 3252 7924 3253 7988
rect 3187 7923 3253 7924
rect 2819 5268 2885 5269
rect 2819 5204 2820 5268
rect 2884 5204 2885 5268
rect 2819 5203 2885 5204
rect 3190 3637 3250 7923
rect 4110 6901 4170 15267
rect 4107 6900 4173 6901
rect 4107 6836 4108 6900
rect 4172 6836 4173 6900
rect 4107 6835 4173 6836
rect 5214 4181 5274 17035
rect 5705 16896 6025 17920
rect 5705 16832 5713 16896
rect 5777 16832 5793 16896
rect 5857 16832 5873 16896
rect 5937 16832 5953 16896
rect 6017 16832 6025 16896
rect 5705 15808 6025 16832
rect 5705 15744 5713 15808
rect 5777 15744 5793 15808
rect 5857 15744 5873 15808
rect 5937 15744 5953 15808
rect 6017 15744 6025 15808
rect 5705 14720 6025 15744
rect 5705 14656 5713 14720
rect 5777 14656 5793 14720
rect 5857 14656 5873 14720
rect 5937 14656 5953 14720
rect 6017 14656 6025 14720
rect 5705 13632 6025 14656
rect 5705 13568 5713 13632
rect 5777 13568 5793 13632
rect 5857 13568 5873 13632
rect 5937 13568 5953 13632
rect 6017 13568 6025 13632
rect 5395 12612 5461 12613
rect 5395 12548 5396 12612
rect 5460 12548 5461 12612
rect 5395 12547 5461 12548
rect 5211 4180 5277 4181
rect 5211 4116 5212 4180
rect 5276 4116 5277 4180
rect 5211 4115 5277 4116
rect 3187 3636 3253 3637
rect 3187 3572 3188 3636
rect 3252 3572 3253 3636
rect 3187 3571 3253 3572
rect 5398 2549 5458 12547
rect 5705 12544 6025 13568
rect 5705 12480 5713 12544
rect 5777 12480 5793 12544
rect 5857 12480 5873 12544
rect 5937 12480 5953 12544
rect 6017 12480 6025 12544
rect 5705 11456 6025 12480
rect 5705 11392 5713 11456
rect 5777 11392 5793 11456
rect 5857 11392 5873 11456
rect 5937 11392 5953 11456
rect 6017 11392 6025 11456
rect 5705 10368 6025 11392
rect 5705 10304 5713 10368
rect 5777 10304 5793 10368
rect 5857 10304 5873 10368
rect 5937 10304 5953 10368
rect 6017 10304 6025 10368
rect 5705 9280 6025 10304
rect 5705 9216 5713 9280
rect 5777 9216 5793 9280
rect 5857 9216 5873 9280
rect 5937 9216 5953 9280
rect 6017 9216 6025 9280
rect 5705 8192 6025 9216
rect 5705 8128 5713 8192
rect 5777 8128 5793 8192
rect 5857 8128 5873 8192
rect 5937 8128 5953 8192
rect 6017 8128 6025 8192
rect 5705 7104 6025 8128
rect 5705 7040 5713 7104
rect 5777 7040 5793 7104
rect 5857 7040 5873 7104
rect 5937 7040 5953 7104
rect 6017 7040 6025 7104
rect 5705 6016 6025 7040
rect 5705 5952 5713 6016
rect 5777 5952 5793 6016
rect 5857 5952 5873 6016
rect 5937 5952 5953 6016
rect 6017 5952 6025 6016
rect 5705 4928 6025 5952
rect 6318 5405 6378 26283
rect 10466 26144 10786 26704
rect 15227 26688 15547 26704
rect 15227 26624 15235 26688
rect 15299 26624 15315 26688
rect 15379 26624 15395 26688
rect 15459 26624 15475 26688
rect 15539 26624 15547 26688
rect 12019 26484 12085 26485
rect 12019 26420 12020 26484
rect 12084 26420 12085 26484
rect 12019 26419 12085 26420
rect 10466 26080 10474 26144
rect 10538 26080 10554 26144
rect 10618 26080 10634 26144
rect 10698 26080 10714 26144
rect 10778 26080 10786 26144
rect 10466 25056 10786 26080
rect 10466 24992 10474 25056
rect 10538 24992 10554 25056
rect 10618 24992 10634 25056
rect 10698 24992 10714 25056
rect 10778 24992 10786 25056
rect 10466 23968 10786 24992
rect 10466 23904 10474 23968
rect 10538 23904 10554 23968
rect 10618 23904 10634 23968
rect 10698 23904 10714 23968
rect 10778 23904 10786 23968
rect 10466 22880 10786 23904
rect 10466 22816 10474 22880
rect 10538 22816 10554 22880
rect 10618 22816 10634 22880
rect 10698 22816 10714 22880
rect 10778 22816 10786 22880
rect 10466 21792 10786 22816
rect 10466 21728 10474 21792
rect 10538 21728 10554 21792
rect 10618 21728 10634 21792
rect 10698 21728 10714 21792
rect 10778 21728 10786 21792
rect 10466 20704 10786 21728
rect 10466 20640 10474 20704
rect 10538 20640 10554 20704
rect 10618 20640 10634 20704
rect 10698 20640 10714 20704
rect 10778 20640 10786 20704
rect 10466 19616 10786 20640
rect 10466 19552 10474 19616
rect 10538 19552 10554 19616
rect 10618 19552 10634 19616
rect 10698 19552 10714 19616
rect 10778 19552 10786 19616
rect 10466 18528 10786 19552
rect 10466 18464 10474 18528
rect 10538 18464 10554 18528
rect 10618 18464 10634 18528
rect 10698 18464 10714 18528
rect 10778 18464 10786 18528
rect 10466 17440 10786 18464
rect 10466 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10786 17440
rect 6499 17236 6565 17237
rect 6499 17172 6500 17236
rect 6564 17172 6565 17236
rect 6499 17171 6565 17172
rect 6502 6765 6562 17171
rect 10466 16352 10786 17376
rect 10466 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10786 16352
rect 10466 15264 10786 16288
rect 10466 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10786 15264
rect 10466 14176 10786 15200
rect 10466 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10786 14176
rect 10466 13088 10786 14112
rect 10466 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10786 13088
rect 8891 12748 8957 12749
rect 8891 12684 8892 12748
rect 8956 12684 8957 12748
rect 8891 12683 8957 12684
rect 7603 11252 7669 11253
rect 7603 11188 7604 11252
rect 7668 11188 7669 11252
rect 7603 11187 7669 11188
rect 7051 8668 7117 8669
rect 7051 8604 7052 8668
rect 7116 8604 7117 8668
rect 7051 8603 7117 8604
rect 7054 6765 7114 8603
rect 6499 6764 6565 6765
rect 6499 6700 6500 6764
rect 6564 6700 6565 6764
rect 6499 6699 6565 6700
rect 7051 6764 7117 6765
rect 7051 6700 7052 6764
rect 7116 6700 7117 6764
rect 7051 6699 7117 6700
rect 6315 5404 6381 5405
rect 6315 5340 6316 5404
rect 6380 5340 6381 5404
rect 6315 5339 6381 5340
rect 7606 4997 7666 11187
rect 8894 5677 8954 12683
rect 9443 12068 9509 12069
rect 9443 12004 9444 12068
rect 9508 12004 9509 12068
rect 9443 12003 9509 12004
rect 9446 8261 9506 12003
rect 10466 12000 10786 13024
rect 10466 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10786 12000
rect 9627 11932 9693 11933
rect 9627 11868 9628 11932
rect 9692 11868 9693 11932
rect 9627 11867 9693 11868
rect 9443 8260 9509 8261
rect 9443 8196 9444 8260
rect 9508 8196 9509 8260
rect 9443 8195 9509 8196
rect 9630 6765 9690 11867
rect 9811 11388 9877 11389
rect 9811 11324 9812 11388
rect 9876 11324 9877 11388
rect 9811 11323 9877 11324
rect 9814 9893 9874 11323
rect 9995 11252 10061 11253
rect 9995 11188 9996 11252
rect 10060 11188 10061 11252
rect 9995 11187 10061 11188
rect 9811 9892 9877 9893
rect 9811 9828 9812 9892
rect 9876 9828 9877 9892
rect 9811 9827 9877 9828
rect 9998 9757 10058 11187
rect 10179 11116 10245 11117
rect 10179 11052 10180 11116
rect 10244 11052 10245 11116
rect 10179 11051 10245 11052
rect 9995 9756 10061 9757
rect 9995 9692 9996 9756
rect 10060 9692 10061 9756
rect 9995 9691 10061 9692
rect 9627 6764 9693 6765
rect 9627 6700 9628 6764
rect 9692 6700 9693 6764
rect 9627 6699 9693 6700
rect 9630 5677 9690 6699
rect 8891 5676 8957 5677
rect 8891 5612 8892 5676
rect 8956 5612 8957 5676
rect 8891 5611 8957 5612
rect 9627 5676 9693 5677
rect 9627 5612 9628 5676
rect 9692 5612 9693 5676
rect 9627 5611 9693 5612
rect 7603 4996 7669 4997
rect 7603 4932 7604 4996
rect 7668 4932 7669 4996
rect 7603 4931 7669 4932
rect 5705 4864 5713 4928
rect 5777 4864 5793 4928
rect 5857 4864 5873 4928
rect 5937 4864 5953 4928
rect 6017 4864 6025 4928
rect 5705 3840 6025 4864
rect 5705 3776 5713 3840
rect 5777 3776 5793 3840
rect 5857 3776 5873 3840
rect 5937 3776 5953 3840
rect 6017 3776 6025 3840
rect 5705 2752 6025 3776
rect 5705 2688 5713 2752
rect 5777 2688 5793 2752
rect 5857 2688 5873 2752
rect 5937 2688 5953 2752
rect 6017 2688 6025 2752
rect 5395 2548 5461 2549
rect 5395 2484 5396 2548
rect 5460 2484 5461 2548
rect 5395 2483 5461 2484
rect 5705 2128 6025 2688
rect 10182 1869 10242 11051
rect 10466 10912 10786 11936
rect 11099 11524 11165 11525
rect 11099 11460 11100 11524
rect 11164 11460 11165 11524
rect 11099 11459 11165 11460
rect 10466 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10786 10912
rect 10466 9824 10786 10848
rect 10466 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10786 9824
rect 10466 8736 10786 9760
rect 10466 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10786 8736
rect 10466 7648 10786 8672
rect 10466 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10786 7648
rect 10466 6560 10786 7584
rect 10466 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10786 6560
rect 10466 5472 10786 6496
rect 11102 5677 11162 11459
rect 12022 10981 12082 26419
rect 14779 26348 14845 26349
rect 14779 26284 14780 26348
rect 14844 26284 14845 26348
rect 14779 26283 14845 26284
rect 13123 24716 13189 24717
rect 13123 24652 13124 24716
rect 13188 24652 13189 24716
rect 13123 24651 13189 24652
rect 12755 20908 12821 20909
rect 12755 20844 12756 20908
rect 12820 20844 12821 20908
rect 12755 20843 12821 20844
rect 12203 16692 12269 16693
rect 12203 16628 12204 16692
rect 12268 16628 12269 16692
rect 12203 16627 12269 16628
rect 12019 10980 12085 10981
rect 12019 10916 12020 10980
rect 12084 10916 12085 10980
rect 12019 10915 12085 10916
rect 12019 9892 12085 9893
rect 12019 9828 12020 9892
rect 12084 9828 12085 9892
rect 12019 9827 12085 9828
rect 11099 5676 11165 5677
rect 11099 5612 11100 5676
rect 11164 5612 11165 5676
rect 11099 5611 11165 5612
rect 10466 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10786 5472
rect 10466 4384 10786 5408
rect 10466 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10786 4384
rect 10466 3296 10786 4320
rect 12022 3909 12082 9827
rect 12206 4045 12266 16627
rect 12571 13972 12637 13973
rect 12571 13908 12572 13972
rect 12636 13908 12637 13972
rect 12571 13907 12637 13908
rect 12574 12610 12634 13907
rect 12390 12550 12634 12610
rect 12390 12450 12450 12550
rect 12390 12390 12634 12450
rect 12574 7037 12634 12390
rect 12758 9621 12818 20843
rect 12939 15060 13005 15061
rect 12939 14996 12940 15060
rect 13004 14996 13005 15060
rect 12939 14995 13005 14996
rect 12942 10845 13002 14995
rect 12939 10844 13005 10845
rect 12939 10780 12940 10844
rect 13004 10780 13005 10844
rect 12939 10779 13005 10780
rect 13126 9621 13186 24651
rect 13307 19276 13373 19277
rect 13307 19212 13308 19276
rect 13372 19212 13373 19276
rect 13307 19211 13373 19212
rect 14411 19276 14477 19277
rect 14411 19212 14412 19276
rect 14476 19212 14477 19276
rect 14411 19211 14477 19212
rect 12755 9620 12821 9621
rect 12755 9556 12756 9620
rect 12820 9556 12821 9620
rect 12755 9555 12821 9556
rect 13123 9620 13189 9621
rect 13123 9556 13124 9620
rect 13188 9556 13189 9620
rect 13123 9555 13189 9556
rect 12571 7036 12637 7037
rect 12571 6972 12572 7036
rect 12636 6972 12637 7036
rect 12571 6971 12637 6972
rect 13310 5405 13370 19211
rect 13859 12068 13925 12069
rect 13859 12004 13860 12068
rect 13924 12004 13925 12068
rect 13859 12003 13925 12004
rect 13491 9484 13557 9485
rect 13491 9420 13492 9484
rect 13556 9420 13557 9484
rect 13491 9419 13557 9420
rect 13494 8125 13554 9419
rect 13491 8124 13557 8125
rect 13491 8060 13492 8124
rect 13556 8060 13557 8124
rect 13491 8059 13557 8060
rect 13862 6493 13922 12003
rect 14414 10845 14474 19211
rect 14595 13972 14661 13973
rect 14595 13908 14596 13972
rect 14660 13908 14661 13972
rect 14595 13907 14661 13908
rect 14598 12341 14658 13907
rect 14782 13565 14842 26283
rect 15227 25600 15547 26624
rect 18643 26348 18709 26349
rect 18643 26284 18644 26348
rect 18708 26284 18709 26348
rect 18643 26283 18709 26284
rect 15227 25536 15235 25600
rect 15299 25536 15315 25600
rect 15379 25536 15395 25600
rect 15459 25536 15475 25600
rect 15539 25536 15547 25600
rect 15227 24512 15547 25536
rect 16619 24716 16685 24717
rect 16619 24652 16620 24716
rect 16684 24652 16685 24716
rect 16619 24651 16685 24652
rect 15227 24448 15235 24512
rect 15299 24448 15315 24512
rect 15379 24448 15395 24512
rect 15459 24448 15475 24512
rect 15539 24448 15547 24512
rect 15227 23424 15547 24448
rect 15227 23360 15235 23424
rect 15299 23360 15315 23424
rect 15379 23360 15395 23424
rect 15459 23360 15475 23424
rect 15539 23360 15547 23424
rect 15227 22336 15547 23360
rect 15227 22272 15235 22336
rect 15299 22272 15315 22336
rect 15379 22272 15395 22336
rect 15459 22272 15475 22336
rect 15539 22272 15547 22336
rect 15227 21248 15547 22272
rect 15227 21184 15235 21248
rect 15299 21184 15315 21248
rect 15379 21184 15395 21248
rect 15459 21184 15475 21248
rect 15539 21184 15547 21248
rect 15227 20160 15547 21184
rect 15227 20096 15235 20160
rect 15299 20096 15315 20160
rect 15379 20096 15395 20160
rect 15459 20096 15475 20160
rect 15539 20096 15547 20160
rect 14963 19684 15029 19685
rect 14963 19620 14964 19684
rect 15028 19620 15029 19684
rect 14963 19619 15029 19620
rect 14779 13564 14845 13565
rect 14779 13500 14780 13564
rect 14844 13500 14845 13564
rect 14779 13499 14845 13500
rect 14595 12340 14661 12341
rect 14595 12276 14596 12340
rect 14660 12276 14661 12340
rect 14595 12275 14661 12276
rect 14411 10844 14477 10845
rect 14411 10780 14412 10844
rect 14476 10780 14477 10844
rect 14411 10779 14477 10780
rect 14043 9348 14109 9349
rect 14043 9284 14044 9348
rect 14108 9284 14109 9348
rect 14043 9283 14109 9284
rect 13859 6492 13925 6493
rect 13859 6428 13860 6492
rect 13924 6428 13925 6492
rect 13859 6427 13925 6428
rect 13307 5404 13373 5405
rect 13307 5340 13308 5404
rect 13372 5340 13373 5404
rect 13307 5339 13373 5340
rect 13310 4861 13370 5339
rect 13307 4860 13373 4861
rect 13307 4796 13308 4860
rect 13372 4796 13373 4860
rect 13307 4795 13373 4796
rect 12203 4044 12269 4045
rect 12203 3980 12204 4044
rect 12268 3980 12269 4044
rect 12203 3979 12269 3980
rect 12019 3908 12085 3909
rect 12019 3844 12020 3908
rect 12084 3844 12085 3908
rect 12019 3843 12085 3844
rect 10466 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10786 3296
rect 10466 2208 10786 3232
rect 14046 3093 14106 9283
rect 14966 9210 15026 19619
rect 15227 19072 15547 20096
rect 15227 19008 15235 19072
rect 15299 19008 15315 19072
rect 15379 19008 15395 19072
rect 15459 19008 15475 19072
rect 15539 19008 15547 19072
rect 15227 17984 15547 19008
rect 15883 18868 15949 18869
rect 15883 18804 15884 18868
rect 15948 18804 15949 18868
rect 15883 18803 15949 18804
rect 15227 17920 15235 17984
rect 15299 17920 15315 17984
rect 15379 17920 15395 17984
rect 15459 17920 15475 17984
rect 15539 17920 15547 17984
rect 15227 16896 15547 17920
rect 15227 16832 15235 16896
rect 15299 16832 15315 16896
rect 15379 16832 15395 16896
rect 15459 16832 15475 16896
rect 15539 16832 15547 16896
rect 15227 15808 15547 16832
rect 15227 15744 15235 15808
rect 15299 15744 15315 15808
rect 15379 15744 15395 15808
rect 15459 15744 15475 15808
rect 15539 15744 15547 15808
rect 15227 14720 15547 15744
rect 15227 14656 15235 14720
rect 15299 14656 15315 14720
rect 15379 14656 15395 14720
rect 15459 14656 15475 14720
rect 15539 14656 15547 14720
rect 15227 13632 15547 14656
rect 15227 13568 15235 13632
rect 15299 13568 15315 13632
rect 15379 13568 15395 13632
rect 15459 13568 15475 13632
rect 15539 13568 15547 13632
rect 15227 12544 15547 13568
rect 15699 13564 15765 13565
rect 15699 13500 15700 13564
rect 15764 13500 15765 13564
rect 15699 13499 15765 13500
rect 15702 13021 15762 13499
rect 15699 13020 15765 13021
rect 15699 12956 15700 13020
rect 15764 12956 15765 13020
rect 15699 12955 15765 12956
rect 15699 12612 15765 12613
rect 15699 12548 15700 12612
rect 15764 12548 15765 12612
rect 15699 12547 15765 12548
rect 15227 12480 15235 12544
rect 15299 12480 15315 12544
rect 15379 12480 15395 12544
rect 15459 12480 15475 12544
rect 15539 12480 15547 12544
rect 15227 11456 15547 12480
rect 15227 11392 15235 11456
rect 15299 11392 15315 11456
rect 15379 11392 15395 11456
rect 15459 11392 15475 11456
rect 15539 11392 15547 11456
rect 15227 10368 15547 11392
rect 15702 10845 15762 12547
rect 15699 10844 15765 10845
rect 15699 10780 15700 10844
rect 15764 10780 15765 10844
rect 15699 10779 15765 10780
rect 15227 10304 15235 10368
rect 15299 10304 15315 10368
rect 15379 10304 15395 10368
rect 15459 10304 15475 10368
rect 15539 10304 15547 10368
rect 15227 9280 15547 10304
rect 15699 9620 15765 9621
rect 15699 9556 15700 9620
rect 15764 9556 15765 9620
rect 15699 9555 15765 9556
rect 15227 9216 15235 9280
rect 15299 9216 15315 9280
rect 15379 9216 15395 9280
rect 15459 9216 15475 9280
rect 15539 9216 15547 9280
rect 14966 9150 15164 9210
rect 15104 9077 15164 9150
rect 15101 9076 15167 9077
rect 15101 9012 15102 9076
rect 15166 9012 15167 9076
rect 15101 9011 15167 9012
rect 15227 8192 15547 9216
rect 15227 8128 15235 8192
rect 15299 8128 15315 8192
rect 15379 8128 15395 8192
rect 15459 8128 15475 8192
rect 15539 8128 15547 8192
rect 15227 7104 15547 8128
rect 15227 7040 15235 7104
rect 15299 7040 15315 7104
rect 15379 7040 15395 7104
rect 15459 7040 15475 7104
rect 15539 7040 15547 7104
rect 15227 6016 15547 7040
rect 15702 6765 15762 9555
rect 15699 6764 15765 6765
rect 15699 6700 15700 6764
rect 15764 6700 15765 6764
rect 15699 6699 15765 6700
rect 15227 5952 15235 6016
rect 15299 5952 15315 6016
rect 15379 5952 15395 6016
rect 15459 5952 15475 6016
rect 15539 5952 15547 6016
rect 15227 4928 15547 5952
rect 15886 5541 15946 18803
rect 16067 18732 16133 18733
rect 16067 18668 16068 18732
rect 16132 18668 16133 18732
rect 16067 18667 16133 18668
rect 16070 11117 16130 18667
rect 16435 15196 16501 15197
rect 16435 15132 16436 15196
rect 16500 15132 16501 15196
rect 16435 15131 16501 15132
rect 16438 12341 16498 15131
rect 16435 12340 16501 12341
rect 16435 12276 16436 12340
rect 16500 12276 16501 12340
rect 16435 12275 16501 12276
rect 16067 11116 16133 11117
rect 16067 11052 16068 11116
rect 16132 11052 16133 11116
rect 16067 11051 16133 11052
rect 16622 5541 16682 24651
rect 17171 24172 17237 24173
rect 17171 24108 17172 24172
rect 17236 24108 17237 24172
rect 17171 24107 17237 24108
rect 16987 18188 17053 18189
rect 16987 18124 16988 18188
rect 17052 18124 17053 18188
rect 16987 18123 17053 18124
rect 16803 13700 16869 13701
rect 16803 13636 16804 13700
rect 16868 13636 16869 13700
rect 16803 13635 16869 13636
rect 16806 11117 16866 13635
rect 16990 11117 17050 18123
rect 16803 11116 16869 11117
rect 16803 11052 16804 11116
rect 16868 11052 16869 11116
rect 16803 11051 16869 11052
rect 16987 11116 17053 11117
rect 16987 11052 16988 11116
rect 17052 11052 17053 11116
rect 16987 11051 17053 11052
rect 15883 5540 15949 5541
rect 15883 5476 15884 5540
rect 15948 5476 15949 5540
rect 15883 5475 15949 5476
rect 16619 5540 16685 5541
rect 16619 5476 16620 5540
rect 16684 5476 16685 5540
rect 16619 5475 16685 5476
rect 15227 4864 15235 4928
rect 15299 4864 15315 4928
rect 15379 4864 15395 4928
rect 15459 4864 15475 4928
rect 15539 4864 15547 4928
rect 15227 3840 15547 4864
rect 15227 3776 15235 3840
rect 15299 3776 15315 3840
rect 15379 3776 15395 3840
rect 15459 3776 15475 3840
rect 15539 3776 15547 3840
rect 14043 3092 14109 3093
rect 14043 3028 14044 3092
rect 14108 3028 14109 3092
rect 14043 3027 14109 3028
rect 10466 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10786 2208
rect 10466 2128 10786 2144
rect 15227 2752 15547 3776
rect 15227 2688 15235 2752
rect 15299 2688 15315 2752
rect 15379 2688 15395 2752
rect 15459 2688 15475 2752
rect 15539 2688 15547 2752
rect 15227 2128 15547 2688
rect 17174 2685 17234 24107
rect 17907 20772 17973 20773
rect 17907 20708 17908 20772
rect 17972 20708 17973 20772
rect 17907 20707 17973 20708
rect 17723 18188 17789 18189
rect 17723 18124 17724 18188
rect 17788 18124 17789 18188
rect 17723 18123 17789 18124
rect 17726 12069 17786 18123
rect 17723 12068 17789 12069
rect 17723 12004 17724 12068
rect 17788 12004 17789 12068
rect 17723 12003 17789 12004
rect 17910 4045 17970 20707
rect 18275 17780 18341 17781
rect 18275 17716 18276 17780
rect 18340 17716 18341 17780
rect 18275 17715 18341 17716
rect 18278 4045 18338 17715
rect 18646 8941 18706 26283
rect 19988 26144 20308 26704
rect 19988 26080 19996 26144
rect 20060 26080 20076 26144
rect 20140 26080 20156 26144
rect 20220 26080 20236 26144
rect 20300 26080 20308 26144
rect 19988 25056 20308 26080
rect 24749 26688 25069 26704
rect 24749 26624 24757 26688
rect 24821 26624 24837 26688
rect 24901 26624 24917 26688
rect 24981 26624 24997 26688
rect 25061 26624 25069 26688
rect 24749 25600 25069 26624
rect 24749 25536 24757 25600
rect 24821 25536 24837 25600
rect 24901 25536 24917 25600
rect 24981 25536 24997 25600
rect 25061 25536 25069 25600
rect 23979 25260 24045 25261
rect 23979 25196 23980 25260
rect 24044 25196 24045 25260
rect 23979 25195 24045 25196
rect 19988 24992 19996 25056
rect 20060 24992 20076 25056
rect 20140 24992 20156 25056
rect 20220 24992 20236 25056
rect 20300 24992 20308 25056
rect 19988 23968 20308 24992
rect 19988 23904 19996 23968
rect 20060 23904 20076 23968
rect 20140 23904 20156 23968
rect 20220 23904 20236 23968
rect 20300 23904 20308 23968
rect 18827 23492 18893 23493
rect 18827 23428 18828 23492
rect 18892 23428 18893 23492
rect 18827 23427 18893 23428
rect 18830 13565 18890 23427
rect 19988 22880 20308 23904
rect 19988 22816 19996 22880
rect 20060 22816 20076 22880
rect 20140 22816 20156 22880
rect 20220 22816 20236 22880
rect 20300 22816 20308 22880
rect 19988 21792 20308 22816
rect 19988 21728 19996 21792
rect 20060 21728 20076 21792
rect 20140 21728 20156 21792
rect 20220 21728 20236 21792
rect 20300 21728 20308 21792
rect 19988 20704 20308 21728
rect 22691 21044 22757 21045
rect 22691 20980 22692 21044
rect 22756 20980 22757 21044
rect 22691 20979 22757 20980
rect 19988 20640 19996 20704
rect 20060 20640 20076 20704
rect 20140 20640 20156 20704
rect 20220 20640 20236 20704
rect 20300 20640 20308 20704
rect 19988 19616 20308 20640
rect 19988 19552 19996 19616
rect 20060 19552 20076 19616
rect 20140 19552 20156 19616
rect 20220 19552 20236 19616
rect 20300 19552 20308 19616
rect 19988 18528 20308 19552
rect 19988 18464 19996 18528
rect 20060 18464 20076 18528
rect 20140 18464 20156 18528
rect 20220 18464 20236 18528
rect 20300 18464 20308 18528
rect 19988 17440 20308 18464
rect 22323 18324 22389 18325
rect 22323 18260 22324 18324
rect 22388 18260 22389 18324
rect 22323 18259 22389 18260
rect 19988 17376 19996 17440
rect 20060 17376 20076 17440
rect 20140 17376 20156 17440
rect 20220 17376 20236 17440
rect 20300 17376 20308 17440
rect 19563 17372 19629 17373
rect 19563 17308 19564 17372
rect 19628 17308 19629 17372
rect 19563 17307 19629 17308
rect 19379 16692 19445 16693
rect 19379 16628 19380 16692
rect 19444 16628 19445 16692
rect 19379 16627 19445 16628
rect 19382 15197 19442 16627
rect 19379 15196 19445 15197
rect 19379 15132 19380 15196
rect 19444 15132 19445 15196
rect 19379 15131 19445 15132
rect 19566 15061 19626 17307
rect 19988 16352 20308 17376
rect 19988 16288 19996 16352
rect 20060 16288 20076 16352
rect 20140 16288 20156 16352
rect 20220 16288 20236 16352
rect 20300 16288 20308 16352
rect 19988 15264 20308 16288
rect 19988 15200 19996 15264
rect 20060 15200 20076 15264
rect 20140 15200 20156 15264
rect 20220 15200 20236 15264
rect 20300 15200 20308 15264
rect 19563 15060 19629 15061
rect 19563 14996 19564 15060
rect 19628 14996 19629 15060
rect 19563 14995 19629 14996
rect 19988 14176 20308 15200
rect 20667 14788 20733 14789
rect 20667 14724 20668 14788
rect 20732 14724 20733 14788
rect 20667 14723 20733 14724
rect 19988 14112 19996 14176
rect 20060 14112 20076 14176
rect 20140 14112 20156 14176
rect 20220 14112 20236 14176
rect 20300 14112 20308 14176
rect 18827 13564 18893 13565
rect 18827 13500 18828 13564
rect 18892 13500 18893 13564
rect 18827 13499 18893 13500
rect 19988 13088 20308 14112
rect 19988 13024 19996 13088
rect 20060 13024 20076 13088
rect 20140 13024 20156 13088
rect 20220 13024 20236 13088
rect 20300 13024 20308 13088
rect 19563 12748 19629 12749
rect 19563 12684 19564 12748
rect 19628 12684 19629 12748
rect 19563 12683 19629 12684
rect 18643 8940 18709 8941
rect 18643 8876 18644 8940
rect 18708 8876 18709 8940
rect 18643 8875 18709 8876
rect 19566 6357 19626 12683
rect 19988 12000 20308 13024
rect 19988 11936 19996 12000
rect 20060 11936 20076 12000
rect 20140 11936 20156 12000
rect 20220 11936 20236 12000
rect 20300 11936 20308 12000
rect 19988 10912 20308 11936
rect 19988 10848 19996 10912
rect 20060 10848 20076 10912
rect 20140 10848 20156 10912
rect 20220 10848 20236 10912
rect 20300 10848 20308 10912
rect 19988 9824 20308 10848
rect 19988 9760 19996 9824
rect 20060 9760 20076 9824
rect 20140 9760 20156 9824
rect 20220 9760 20236 9824
rect 20300 9760 20308 9824
rect 19988 8736 20308 9760
rect 20670 8805 20730 14723
rect 20667 8804 20733 8805
rect 20667 8740 20668 8804
rect 20732 8740 20733 8804
rect 20667 8739 20733 8740
rect 19988 8672 19996 8736
rect 20060 8672 20076 8736
rect 20140 8672 20156 8736
rect 20220 8672 20236 8736
rect 20300 8672 20308 8736
rect 19988 7648 20308 8672
rect 19988 7584 19996 7648
rect 20060 7584 20076 7648
rect 20140 7584 20156 7648
rect 20220 7584 20236 7648
rect 20300 7584 20308 7648
rect 19988 6560 20308 7584
rect 22326 6629 22386 18259
rect 22694 9621 22754 20979
rect 23427 12204 23493 12205
rect 23427 12140 23428 12204
rect 23492 12140 23493 12204
rect 23427 12139 23493 12140
rect 22691 9620 22757 9621
rect 22691 9556 22692 9620
rect 22756 9556 22757 9620
rect 22691 9555 22757 9556
rect 23430 7717 23490 12139
rect 23427 7716 23493 7717
rect 23427 7652 23428 7716
rect 23492 7652 23493 7716
rect 23427 7651 23493 7652
rect 22323 6628 22389 6629
rect 22323 6564 22324 6628
rect 22388 6564 22389 6628
rect 22323 6563 22389 6564
rect 19988 6496 19996 6560
rect 20060 6496 20076 6560
rect 20140 6496 20156 6560
rect 20220 6496 20236 6560
rect 20300 6496 20308 6560
rect 19563 6356 19629 6357
rect 19563 6292 19564 6356
rect 19628 6292 19629 6356
rect 19563 6291 19629 6292
rect 19988 5472 20308 6496
rect 19988 5408 19996 5472
rect 20060 5408 20076 5472
rect 20140 5408 20156 5472
rect 20220 5408 20236 5472
rect 20300 5408 20308 5472
rect 19988 4384 20308 5408
rect 19988 4320 19996 4384
rect 20060 4320 20076 4384
rect 20140 4320 20156 4384
rect 20220 4320 20236 4384
rect 20300 4320 20308 4384
rect 17907 4044 17973 4045
rect 17907 3980 17908 4044
rect 17972 3980 17973 4044
rect 17907 3979 17973 3980
rect 18275 4044 18341 4045
rect 18275 3980 18276 4044
rect 18340 3980 18341 4044
rect 18275 3979 18341 3980
rect 19988 3296 20308 4320
rect 19988 3232 19996 3296
rect 20060 3232 20076 3296
rect 20140 3232 20156 3296
rect 20220 3232 20236 3296
rect 20300 3232 20308 3296
rect 17171 2684 17237 2685
rect 17171 2620 17172 2684
rect 17236 2620 17237 2684
rect 17171 2619 17237 2620
rect 19988 2208 20308 3232
rect 23982 2549 24042 25195
rect 24749 24512 25069 25536
rect 24749 24448 24757 24512
rect 24821 24448 24837 24512
rect 24901 24448 24917 24512
rect 24981 24448 24997 24512
rect 25061 24448 25069 24512
rect 24749 23424 25069 24448
rect 24749 23360 24757 23424
rect 24821 23360 24837 23424
rect 24901 23360 24917 23424
rect 24981 23360 24997 23424
rect 25061 23360 25069 23424
rect 24749 22336 25069 23360
rect 29510 26144 29830 26704
rect 29510 26080 29518 26144
rect 29582 26080 29598 26144
rect 29662 26080 29678 26144
rect 29742 26080 29758 26144
rect 29822 26080 29830 26144
rect 29510 25056 29830 26080
rect 29510 24992 29518 25056
rect 29582 24992 29598 25056
rect 29662 24992 29678 25056
rect 29742 24992 29758 25056
rect 29822 24992 29830 25056
rect 29510 23968 29830 24992
rect 29510 23904 29518 23968
rect 29582 23904 29598 23968
rect 29662 23904 29678 23968
rect 29742 23904 29758 23968
rect 29822 23904 29830 23968
rect 25635 22948 25701 22949
rect 25635 22884 25636 22948
rect 25700 22884 25701 22948
rect 25635 22883 25701 22884
rect 24749 22272 24757 22336
rect 24821 22272 24837 22336
rect 24901 22272 24917 22336
rect 24981 22272 24997 22336
rect 25061 22272 25069 22336
rect 24749 21248 25069 22272
rect 24749 21184 24757 21248
rect 24821 21184 24837 21248
rect 24901 21184 24917 21248
rect 24981 21184 24997 21248
rect 25061 21184 25069 21248
rect 24749 20160 25069 21184
rect 24749 20096 24757 20160
rect 24821 20096 24837 20160
rect 24901 20096 24917 20160
rect 24981 20096 24997 20160
rect 25061 20096 25069 20160
rect 24749 19072 25069 20096
rect 24749 19008 24757 19072
rect 24821 19008 24837 19072
rect 24901 19008 24917 19072
rect 24981 19008 24997 19072
rect 25061 19008 25069 19072
rect 24749 17984 25069 19008
rect 25451 18596 25517 18597
rect 25451 18532 25452 18596
rect 25516 18532 25517 18596
rect 25451 18531 25517 18532
rect 24749 17920 24757 17984
rect 24821 17920 24837 17984
rect 24901 17920 24917 17984
rect 24981 17920 24997 17984
rect 25061 17920 25069 17984
rect 24749 16896 25069 17920
rect 24749 16832 24757 16896
rect 24821 16832 24837 16896
rect 24901 16832 24917 16896
rect 24981 16832 24997 16896
rect 25061 16832 25069 16896
rect 24749 15808 25069 16832
rect 24749 15744 24757 15808
rect 24821 15744 24837 15808
rect 24901 15744 24917 15808
rect 24981 15744 24997 15808
rect 25061 15744 25069 15808
rect 24749 14720 25069 15744
rect 24749 14656 24757 14720
rect 24821 14656 24837 14720
rect 24901 14656 24917 14720
rect 24981 14656 24997 14720
rect 25061 14656 25069 14720
rect 24749 13632 25069 14656
rect 24749 13568 24757 13632
rect 24821 13568 24837 13632
rect 24901 13568 24917 13632
rect 24981 13568 24997 13632
rect 25061 13568 25069 13632
rect 24749 12544 25069 13568
rect 24749 12480 24757 12544
rect 24821 12480 24837 12544
rect 24901 12480 24917 12544
rect 24981 12480 24997 12544
rect 25061 12480 25069 12544
rect 24749 11456 25069 12480
rect 24749 11392 24757 11456
rect 24821 11392 24837 11456
rect 24901 11392 24917 11456
rect 24981 11392 24997 11456
rect 25061 11392 25069 11456
rect 24749 10368 25069 11392
rect 25454 10981 25514 18531
rect 25451 10980 25517 10981
rect 25451 10916 25452 10980
rect 25516 10916 25517 10980
rect 25451 10915 25517 10916
rect 24749 10304 24757 10368
rect 24821 10304 24837 10368
rect 24901 10304 24917 10368
rect 24981 10304 24997 10368
rect 25061 10304 25069 10368
rect 24749 9280 25069 10304
rect 24749 9216 24757 9280
rect 24821 9216 24837 9280
rect 24901 9216 24917 9280
rect 24981 9216 24997 9280
rect 25061 9216 25069 9280
rect 24531 8940 24597 8941
rect 24531 8876 24532 8940
rect 24596 8876 24597 8940
rect 24531 8875 24597 8876
rect 24534 7989 24594 8875
rect 24749 8192 25069 9216
rect 24749 8128 24757 8192
rect 24821 8128 24837 8192
rect 24901 8128 24917 8192
rect 24981 8128 24997 8192
rect 25061 8128 25069 8192
rect 24531 7988 24597 7989
rect 24531 7924 24532 7988
rect 24596 7924 24597 7988
rect 24531 7923 24597 7924
rect 24749 7104 25069 8128
rect 24749 7040 24757 7104
rect 24821 7040 24837 7104
rect 24901 7040 24917 7104
rect 24981 7040 24997 7104
rect 25061 7040 25069 7104
rect 24749 6016 25069 7040
rect 24749 5952 24757 6016
rect 24821 5952 24837 6016
rect 24901 5952 24917 6016
rect 24981 5952 24997 6016
rect 25061 5952 25069 6016
rect 24749 4928 25069 5952
rect 25638 5949 25698 22883
rect 29510 22880 29830 23904
rect 29510 22816 29518 22880
rect 29582 22816 29598 22880
rect 29662 22816 29678 22880
rect 29742 22816 29758 22880
rect 29822 22816 29830 22880
rect 29510 21792 29830 22816
rect 34271 26688 34591 26704
rect 34271 26624 34279 26688
rect 34343 26624 34359 26688
rect 34423 26624 34439 26688
rect 34503 26624 34519 26688
rect 34583 26624 34591 26688
rect 34271 25600 34591 26624
rect 34271 25536 34279 25600
rect 34343 25536 34359 25600
rect 34423 25536 34439 25600
rect 34503 25536 34519 25600
rect 34583 25536 34591 25600
rect 34271 24512 34591 25536
rect 34271 24448 34279 24512
rect 34343 24448 34359 24512
rect 34423 24448 34439 24512
rect 34503 24448 34519 24512
rect 34583 24448 34591 24512
rect 34271 23424 34591 24448
rect 34271 23360 34279 23424
rect 34343 23360 34359 23424
rect 34423 23360 34439 23424
rect 34503 23360 34519 23424
rect 34583 23360 34591 23424
rect 30235 22404 30301 22405
rect 30235 22340 30236 22404
rect 30300 22340 30301 22404
rect 30235 22339 30301 22340
rect 29510 21728 29518 21792
rect 29582 21728 29598 21792
rect 29662 21728 29678 21792
rect 29742 21728 29758 21792
rect 29822 21728 29830 21792
rect 29510 20704 29830 21728
rect 29510 20640 29518 20704
rect 29582 20640 29598 20704
rect 29662 20640 29678 20704
rect 29742 20640 29758 20704
rect 29822 20640 29830 20704
rect 29510 19616 29830 20640
rect 29510 19552 29518 19616
rect 29582 19552 29598 19616
rect 29662 19552 29678 19616
rect 29742 19552 29758 19616
rect 29822 19552 29830 19616
rect 29510 18528 29830 19552
rect 29510 18464 29518 18528
rect 29582 18464 29598 18528
rect 29662 18464 29678 18528
rect 29742 18464 29758 18528
rect 29822 18464 29830 18528
rect 27659 18052 27725 18053
rect 27659 17988 27660 18052
rect 27724 17988 27725 18052
rect 27659 17987 27725 17988
rect 27107 17916 27173 17917
rect 27107 17852 27108 17916
rect 27172 17852 27173 17916
rect 27107 17851 27173 17852
rect 25819 11796 25885 11797
rect 25819 11732 25820 11796
rect 25884 11732 25885 11796
rect 25819 11731 25885 11732
rect 26739 11796 26805 11797
rect 26739 11732 26740 11796
rect 26804 11732 26805 11796
rect 26739 11731 26805 11732
rect 25822 6357 25882 11731
rect 26187 8532 26253 8533
rect 26187 8468 26188 8532
rect 26252 8468 26253 8532
rect 26187 8467 26253 8468
rect 25819 6356 25885 6357
rect 25819 6292 25820 6356
rect 25884 6292 25885 6356
rect 25819 6291 25885 6292
rect 25822 6085 25882 6291
rect 25819 6084 25885 6085
rect 25819 6020 25820 6084
rect 25884 6020 25885 6084
rect 25819 6019 25885 6020
rect 26190 5949 26250 8467
rect 25635 5948 25701 5949
rect 25635 5884 25636 5948
rect 25700 5884 25701 5948
rect 25635 5883 25701 5884
rect 26187 5948 26253 5949
rect 26187 5884 26188 5948
rect 26252 5884 26253 5948
rect 26187 5883 26253 5884
rect 24749 4864 24757 4928
rect 24821 4864 24837 4928
rect 24901 4864 24917 4928
rect 24981 4864 24997 4928
rect 25061 4864 25069 4928
rect 24749 3840 25069 4864
rect 24749 3776 24757 3840
rect 24821 3776 24837 3840
rect 24901 3776 24917 3840
rect 24981 3776 24997 3840
rect 25061 3776 25069 3840
rect 24749 2752 25069 3776
rect 26742 3229 26802 11731
rect 26923 9756 26989 9757
rect 26923 9692 26924 9756
rect 26988 9692 26989 9756
rect 26923 9691 26989 9692
rect 26926 6493 26986 9691
rect 26923 6492 26989 6493
rect 26923 6428 26924 6492
rect 26988 6428 26989 6492
rect 26923 6427 26989 6428
rect 27110 4453 27170 17851
rect 27475 15196 27541 15197
rect 27475 15132 27476 15196
rect 27540 15132 27541 15196
rect 27475 15131 27541 15132
rect 27478 10845 27538 15131
rect 27475 10844 27541 10845
rect 27475 10780 27476 10844
rect 27540 10780 27541 10844
rect 27475 10779 27541 10780
rect 27107 4452 27173 4453
rect 27107 4388 27108 4452
rect 27172 4388 27173 4452
rect 27107 4387 27173 4388
rect 26739 3228 26805 3229
rect 26739 3164 26740 3228
rect 26804 3164 26805 3228
rect 26739 3163 26805 3164
rect 24749 2688 24757 2752
rect 24821 2688 24837 2752
rect 24901 2688 24917 2752
rect 24981 2688 24997 2752
rect 25061 2688 25069 2752
rect 23979 2548 24045 2549
rect 23979 2484 23980 2548
rect 24044 2484 24045 2548
rect 23979 2483 24045 2484
rect 19988 2144 19996 2208
rect 20060 2144 20076 2208
rect 20140 2144 20156 2208
rect 20220 2144 20236 2208
rect 20300 2144 20308 2208
rect 19988 2128 20308 2144
rect 24749 2128 25069 2688
rect 27662 2685 27722 17987
rect 29510 17440 29830 18464
rect 29510 17376 29518 17440
rect 29582 17376 29598 17440
rect 29662 17376 29678 17440
rect 29742 17376 29758 17440
rect 29822 17376 29830 17440
rect 29510 16352 29830 17376
rect 29510 16288 29518 16352
rect 29582 16288 29598 16352
rect 29662 16288 29678 16352
rect 29742 16288 29758 16352
rect 29822 16288 29830 16352
rect 29510 15264 29830 16288
rect 29510 15200 29518 15264
rect 29582 15200 29598 15264
rect 29662 15200 29678 15264
rect 29742 15200 29758 15264
rect 29822 15200 29830 15264
rect 29510 14176 29830 15200
rect 29510 14112 29518 14176
rect 29582 14112 29598 14176
rect 29662 14112 29678 14176
rect 29742 14112 29758 14176
rect 29822 14112 29830 14176
rect 28395 13564 28461 13565
rect 28395 13500 28396 13564
rect 28460 13500 28461 13564
rect 28395 13499 28461 13500
rect 27843 13292 27909 13293
rect 27843 13228 27844 13292
rect 27908 13228 27909 13292
rect 27843 13227 27909 13228
rect 27846 9757 27906 13227
rect 28211 11660 28277 11661
rect 28211 11596 28212 11660
rect 28276 11596 28277 11660
rect 28211 11595 28277 11596
rect 27843 9756 27909 9757
rect 27843 9692 27844 9756
rect 27908 9692 27909 9756
rect 27843 9691 27909 9692
rect 27843 9484 27909 9485
rect 27843 9420 27844 9484
rect 27908 9420 27909 9484
rect 27843 9419 27909 9420
rect 28027 9484 28093 9485
rect 28027 9420 28028 9484
rect 28092 9420 28093 9484
rect 28027 9419 28093 9420
rect 27846 9346 27906 9419
rect 28030 9346 28090 9419
rect 27846 9286 28090 9346
rect 28214 5269 28274 11595
rect 28398 8669 28458 13499
rect 29510 13088 29830 14112
rect 30051 13292 30117 13293
rect 30051 13228 30052 13292
rect 30116 13228 30117 13292
rect 30051 13227 30117 13228
rect 29510 13024 29518 13088
rect 29582 13024 29598 13088
rect 29662 13024 29678 13088
rect 29742 13024 29758 13088
rect 29822 13024 29830 13088
rect 29510 12000 29830 13024
rect 29510 11936 29518 12000
rect 29582 11936 29598 12000
rect 29662 11936 29678 12000
rect 29742 11936 29758 12000
rect 29822 11936 29830 12000
rect 29315 10980 29381 10981
rect 29315 10916 29316 10980
rect 29380 10916 29381 10980
rect 29315 10915 29381 10916
rect 29318 10573 29378 10915
rect 29510 10912 29830 11936
rect 29510 10848 29518 10912
rect 29582 10848 29598 10912
rect 29662 10848 29678 10912
rect 29742 10848 29758 10912
rect 29822 10848 29830 10912
rect 29315 10572 29381 10573
rect 29315 10508 29316 10572
rect 29380 10508 29381 10572
rect 29315 10507 29381 10508
rect 28947 10164 29013 10165
rect 28947 10100 28948 10164
rect 29012 10100 29013 10164
rect 28947 10099 29013 10100
rect 28579 9620 28645 9621
rect 28579 9556 28580 9620
rect 28644 9556 28645 9620
rect 28579 9555 28645 9556
rect 28582 8669 28642 9555
rect 28763 9348 28829 9349
rect 28763 9284 28764 9348
rect 28828 9284 28829 9348
rect 28763 9283 28829 9284
rect 28766 8805 28826 9283
rect 28763 8804 28829 8805
rect 28763 8740 28764 8804
rect 28828 8740 28829 8804
rect 28763 8739 28829 8740
rect 28395 8668 28461 8669
rect 28395 8604 28396 8668
rect 28460 8604 28461 8668
rect 28395 8603 28461 8604
rect 28579 8668 28645 8669
rect 28579 8604 28580 8668
rect 28644 8604 28645 8668
rect 28579 8603 28645 8604
rect 28211 5268 28277 5269
rect 28211 5204 28212 5268
rect 28276 5204 28277 5268
rect 28211 5203 28277 5204
rect 28950 3365 29010 10099
rect 29131 9892 29197 9893
rect 29131 9828 29132 9892
rect 29196 9828 29197 9892
rect 29131 9827 29197 9828
rect 29134 8125 29194 9827
rect 29510 9824 29830 10848
rect 29510 9760 29518 9824
rect 29582 9760 29598 9824
rect 29662 9760 29678 9824
rect 29742 9760 29758 9824
rect 29822 9760 29830 9824
rect 29510 8736 29830 9760
rect 29510 8672 29518 8736
rect 29582 8672 29598 8736
rect 29662 8672 29678 8736
rect 29742 8672 29758 8736
rect 29822 8672 29830 8736
rect 29131 8124 29197 8125
rect 29131 8060 29132 8124
rect 29196 8060 29197 8124
rect 29131 8059 29197 8060
rect 29510 7648 29830 8672
rect 29510 7584 29518 7648
rect 29582 7584 29598 7648
rect 29662 7584 29678 7648
rect 29742 7584 29758 7648
rect 29822 7584 29830 7648
rect 29510 6560 29830 7584
rect 29510 6496 29518 6560
rect 29582 6496 29598 6560
rect 29662 6496 29678 6560
rect 29742 6496 29758 6560
rect 29822 6496 29830 6560
rect 29510 5472 29830 6496
rect 29510 5408 29518 5472
rect 29582 5408 29598 5472
rect 29662 5408 29678 5472
rect 29742 5408 29758 5472
rect 29822 5408 29830 5472
rect 29510 4384 29830 5408
rect 29510 4320 29518 4384
rect 29582 4320 29598 4384
rect 29662 4320 29678 4384
rect 29742 4320 29758 4384
rect 29822 4320 29830 4384
rect 28947 3364 29013 3365
rect 28947 3300 28948 3364
rect 29012 3300 29013 3364
rect 28947 3299 29013 3300
rect 29510 3296 29830 4320
rect 30054 4045 30114 13227
rect 30238 9757 30298 22339
rect 34271 22336 34591 23360
rect 34271 22272 34279 22336
rect 34343 22272 34359 22336
rect 34423 22272 34439 22336
rect 34503 22272 34519 22336
rect 34583 22272 34591 22336
rect 33179 22132 33245 22133
rect 33179 22068 33180 22132
rect 33244 22068 33245 22132
rect 33179 22067 33245 22068
rect 32995 21860 33061 21861
rect 32995 21796 32996 21860
rect 33060 21796 33061 21860
rect 32995 21795 33061 21796
rect 32811 20772 32877 20773
rect 32811 20708 32812 20772
rect 32876 20708 32877 20772
rect 32811 20707 32877 20708
rect 32627 19412 32693 19413
rect 32627 19348 32628 19412
rect 32692 19348 32693 19412
rect 32627 19347 32693 19348
rect 31339 17100 31405 17101
rect 31339 17036 31340 17100
rect 31404 17036 31405 17100
rect 31339 17035 31405 17036
rect 30419 13564 30485 13565
rect 30419 13500 30420 13564
rect 30484 13500 30485 13564
rect 30419 13499 30485 13500
rect 30235 9756 30301 9757
rect 30235 9692 30236 9756
rect 30300 9692 30301 9756
rect 30235 9691 30301 9692
rect 30422 9213 30482 13499
rect 31155 12204 31221 12205
rect 31155 12140 31156 12204
rect 31220 12140 31221 12204
rect 31155 12139 31221 12140
rect 31158 11117 31218 12139
rect 31155 11116 31221 11117
rect 31155 11052 31156 11116
rect 31220 11052 31221 11116
rect 31155 11051 31221 11052
rect 30419 9212 30485 9213
rect 30419 9148 30420 9212
rect 30484 9148 30485 9212
rect 30419 9147 30485 9148
rect 30422 5949 30482 9147
rect 31158 6901 31218 11051
rect 31342 9757 31402 17035
rect 31707 12476 31773 12477
rect 31707 12412 31708 12476
rect 31772 12450 31773 12476
rect 31772 12412 31954 12450
rect 31707 12411 31954 12412
rect 31710 12390 31954 12411
rect 31339 9756 31405 9757
rect 31339 9692 31340 9756
rect 31404 9692 31405 9756
rect 31339 9691 31405 9692
rect 31894 9621 31954 12390
rect 31891 9620 31957 9621
rect 31891 9556 31892 9620
rect 31956 9556 31957 9620
rect 31891 9555 31957 9556
rect 31155 6900 31221 6901
rect 31155 6836 31156 6900
rect 31220 6836 31221 6900
rect 31155 6835 31221 6836
rect 30419 5948 30485 5949
rect 30419 5884 30420 5948
rect 30484 5884 30485 5948
rect 30419 5883 30485 5884
rect 30051 4044 30117 4045
rect 30051 3980 30052 4044
rect 30116 3980 30117 4044
rect 30051 3979 30117 3980
rect 32630 3909 32690 19347
rect 32814 8805 32874 20707
rect 32998 8805 33058 21795
rect 32811 8804 32877 8805
rect 32811 8740 32812 8804
rect 32876 8740 32877 8804
rect 32811 8739 32877 8740
rect 32995 8804 33061 8805
rect 32995 8740 32996 8804
rect 33060 8740 33061 8804
rect 32995 8739 33061 8740
rect 32627 3908 32693 3909
rect 32627 3844 32628 3908
rect 32692 3844 32693 3908
rect 32627 3843 32693 3844
rect 29510 3232 29518 3296
rect 29582 3232 29598 3296
rect 29662 3232 29678 3296
rect 29742 3232 29758 3296
rect 29822 3232 29830 3296
rect 27659 2684 27725 2685
rect 27659 2620 27660 2684
rect 27724 2620 27725 2684
rect 27659 2619 27725 2620
rect 29510 2208 29830 3232
rect 33182 2685 33242 22067
rect 34271 21248 34591 22272
rect 34271 21184 34279 21248
rect 34343 21184 34359 21248
rect 34423 21184 34439 21248
rect 34503 21184 34519 21248
rect 34583 21184 34591 21248
rect 34271 20160 34591 21184
rect 34271 20096 34279 20160
rect 34343 20096 34359 20160
rect 34423 20096 34439 20160
rect 34503 20096 34519 20160
rect 34583 20096 34591 20160
rect 34271 19072 34591 20096
rect 34271 19008 34279 19072
rect 34343 19008 34359 19072
rect 34423 19008 34439 19072
rect 34503 19008 34519 19072
rect 34583 19008 34591 19072
rect 33731 18188 33797 18189
rect 33731 18124 33732 18188
rect 33796 18124 33797 18188
rect 33731 18123 33797 18124
rect 33734 5541 33794 18123
rect 34271 17984 34591 19008
rect 34271 17920 34279 17984
rect 34343 17920 34359 17984
rect 34423 17920 34439 17984
rect 34503 17920 34519 17984
rect 34583 17920 34591 17984
rect 34271 16896 34591 17920
rect 34271 16832 34279 16896
rect 34343 16832 34359 16896
rect 34423 16832 34439 16896
rect 34503 16832 34519 16896
rect 34583 16832 34591 16896
rect 34271 15808 34591 16832
rect 34271 15744 34279 15808
rect 34343 15744 34359 15808
rect 34423 15744 34439 15808
rect 34503 15744 34519 15808
rect 34583 15744 34591 15808
rect 34271 14720 34591 15744
rect 34271 14656 34279 14720
rect 34343 14656 34359 14720
rect 34423 14656 34439 14720
rect 34503 14656 34519 14720
rect 34583 14656 34591 14720
rect 34271 13632 34591 14656
rect 34271 13568 34279 13632
rect 34343 13568 34359 13632
rect 34423 13568 34439 13632
rect 34503 13568 34519 13632
rect 34583 13568 34591 13632
rect 34271 12544 34591 13568
rect 34271 12480 34279 12544
rect 34343 12480 34359 12544
rect 34423 12480 34439 12544
rect 34503 12480 34519 12544
rect 34583 12480 34591 12544
rect 34271 11456 34591 12480
rect 34271 11392 34279 11456
rect 34343 11392 34359 11456
rect 34423 11392 34439 11456
rect 34503 11392 34519 11456
rect 34583 11392 34591 11456
rect 34271 10368 34591 11392
rect 34271 10304 34279 10368
rect 34343 10304 34359 10368
rect 34423 10304 34439 10368
rect 34503 10304 34519 10368
rect 34583 10304 34591 10368
rect 34271 9280 34591 10304
rect 34271 9216 34279 9280
rect 34343 9216 34359 9280
rect 34423 9216 34439 9280
rect 34503 9216 34519 9280
rect 34583 9216 34591 9280
rect 34271 8192 34591 9216
rect 39032 26144 39352 26704
rect 39032 26080 39040 26144
rect 39104 26080 39120 26144
rect 39184 26080 39200 26144
rect 39264 26080 39280 26144
rect 39344 26080 39352 26144
rect 39032 25056 39352 26080
rect 39032 24992 39040 25056
rect 39104 24992 39120 25056
rect 39184 24992 39200 25056
rect 39264 24992 39280 25056
rect 39344 24992 39352 25056
rect 39032 23968 39352 24992
rect 39032 23904 39040 23968
rect 39104 23904 39120 23968
rect 39184 23904 39200 23968
rect 39264 23904 39280 23968
rect 39344 23904 39352 23968
rect 39032 22880 39352 23904
rect 39032 22816 39040 22880
rect 39104 22816 39120 22880
rect 39184 22816 39200 22880
rect 39264 22816 39280 22880
rect 39344 22816 39352 22880
rect 39032 21792 39352 22816
rect 39032 21728 39040 21792
rect 39104 21728 39120 21792
rect 39184 21728 39200 21792
rect 39264 21728 39280 21792
rect 39344 21728 39352 21792
rect 39032 20704 39352 21728
rect 39032 20640 39040 20704
rect 39104 20640 39120 20704
rect 39184 20640 39200 20704
rect 39264 20640 39280 20704
rect 39344 20640 39352 20704
rect 39032 19616 39352 20640
rect 39032 19552 39040 19616
rect 39104 19552 39120 19616
rect 39184 19552 39200 19616
rect 39264 19552 39280 19616
rect 39344 19552 39352 19616
rect 39032 18528 39352 19552
rect 39032 18464 39040 18528
rect 39104 18464 39120 18528
rect 39184 18464 39200 18528
rect 39264 18464 39280 18528
rect 39344 18464 39352 18528
rect 39032 17440 39352 18464
rect 39032 17376 39040 17440
rect 39104 17376 39120 17440
rect 39184 17376 39200 17440
rect 39264 17376 39280 17440
rect 39344 17376 39352 17440
rect 39032 16352 39352 17376
rect 39032 16288 39040 16352
rect 39104 16288 39120 16352
rect 39184 16288 39200 16352
rect 39264 16288 39280 16352
rect 39344 16288 39352 16352
rect 39032 15264 39352 16288
rect 39032 15200 39040 15264
rect 39104 15200 39120 15264
rect 39184 15200 39200 15264
rect 39264 15200 39280 15264
rect 39344 15200 39352 15264
rect 39032 14176 39352 15200
rect 39032 14112 39040 14176
rect 39104 14112 39120 14176
rect 39184 14112 39200 14176
rect 39264 14112 39280 14176
rect 39344 14112 39352 14176
rect 39032 13088 39352 14112
rect 39032 13024 39040 13088
rect 39104 13024 39120 13088
rect 39184 13024 39200 13088
rect 39264 13024 39280 13088
rect 39344 13024 39352 13088
rect 39032 12000 39352 13024
rect 39032 11936 39040 12000
rect 39104 11936 39120 12000
rect 39184 11936 39200 12000
rect 39264 11936 39280 12000
rect 39344 11936 39352 12000
rect 39032 10912 39352 11936
rect 39032 10848 39040 10912
rect 39104 10848 39120 10912
rect 39184 10848 39200 10912
rect 39264 10848 39280 10912
rect 39344 10848 39352 10912
rect 39032 9824 39352 10848
rect 39032 9760 39040 9824
rect 39104 9760 39120 9824
rect 39184 9760 39200 9824
rect 39264 9760 39280 9824
rect 39344 9760 39352 9824
rect 34651 8940 34717 8941
rect 34651 8876 34652 8940
rect 34716 8876 34717 8940
rect 34651 8875 34717 8876
rect 34271 8128 34279 8192
rect 34343 8128 34359 8192
rect 34423 8128 34439 8192
rect 34503 8128 34519 8192
rect 34583 8128 34591 8192
rect 34271 7104 34591 8128
rect 34271 7040 34279 7104
rect 34343 7040 34359 7104
rect 34423 7040 34439 7104
rect 34503 7040 34519 7104
rect 34583 7040 34591 7104
rect 34271 6016 34591 7040
rect 34271 5952 34279 6016
rect 34343 5952 34359 6016
rect 34423 5952 34439 6016
rect 34503 5952 34519 6016
rect 34583 5952 34591 6016
rect 33731 5540 33797 5541
rect 33731 5476 33732 5540
rect 33796 5476 33797 5540
rect 33731 5475 33797 5476
rect 34271 4928 34591 5952
rect 34271 4864 34279 4928
rect 34343 4864 34359 4928
rect 34423 4864 34439 4928
rect 34503 4864 34519 4928
rect 34583 4864 34591 4928
rect 34271 3840 34591 4864
rect 34271 3776 34279 3840
rect 34343 3776 34359 3840
rect 34423 3776 34439 3840
rect 34503 3776 34519 3840
rect 34583 3776 34591 3840
rect 34271 2752 34591 3776
rect 34654 3365 34714 8875
rect 39032 8736 39352 9760
rect 39032 8672 39040 8736
rect 39104 8672 39120 8736
rect 39184 8672 39200 8736
rect 39264 8672 39280 8736
rect 39344 8672 39352 8736
rect 39032 7648 39352 8672
rect 39032 7584 39040 7648
rect 39104 7584 39120 7648
rect 39184 7584 39200 7648
rect 39264 7584 39280 7648
rect 39344 7584 39352 7648
rect 39032 6560 39352 7584
rect 39032 6496 39040 6560
rect 39104 6496 39120 6560
rect 39184 6496 39200 6560
rect 39264 6496 39280 6560
rect 39344 6496 39352 6560
rect 39032 5472 39352 6496
rect 39032 5408 39040 5472
rect 39104 5408 39120 5472
rect 39184 5408 39200 5472
rect 39264 5408 39280 5472
rect 39344 5408 39352 5472
rect 39032 4384 39352 5408
rect 39032 4320 39040 4384
rect 39104 4320 39120 4384
rect 39184 4320 39200 4384
rect 39264 4320 39280 4384
rect 39344 4320 39352 4384
rect 34651 3364 34717 3365
rect 34651 3300 34652 3364
rect 34716 3300 34717 3364
rect 34651 3299 34717 3300
rect 34271 2688 34279 2752
rect 34343 2688 34359 2752
rect 34423 2688 34439 2752
rect 34503 2688 34519 2752
rect 34583 2688 34591 2752
rect 33179 2684 33245 2685
rect 33179 2620 33180 2684
rect 33244 2620 33245 2684
rect 33179 2619 33245 2620
rect 29510 2144 29518 2208
rect 29582 2144 29598 2208
rect 29662 2144 29678 2208
rect 29742 2144 29758 2208
rect 29822 2144 29830 2208
rect 29510 2128 29830 2144
rect 34271 2128 34591 2688
rect 39032 3296 39352 4320
rect 39032 3232 39040 3296
rect 39104 3232 39120 3296
rect 39184 3232 39200 3296
rect 39264 3232 39280 3296
rect 39344 3232 39352 3296
rect 39032 2208 39352 3232
rect 39032 2144 39040 2208
rect 39104 2144 39120 2208
rect 39184 2144 39200 2208
rect 39264 2144 39280 2208
rect 39344 2144 39352 2208
rect 39032 2128 39352 2144
rect 10179 1868 10245 1869
rect 10179 1804 10180 1868
rect 10244 1804 10245 1868
rect 10179 1803 10245 1804
rect 2635 1324 2701 1325
rect 2635 1260 2636 1324
rect 2700 1260 2701 1324
rect 2635 1259 2701 1260
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 36984 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 34684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 28060 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 37996 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 2116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 36064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 5336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 24748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 24748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35
timestamp 1676037725
transform 1 0 4324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43
timestamp 1676037725
transform 1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1676037725
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1676037725
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1676037725
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1676037725
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1676037725
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1676037725
transform 1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_229
timestamp 1676037725
transform 1 0 22172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1676037725
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_303
timestamp 1676037725
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_317
timestamp 1676037725
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_327
timestamp 1676037725
transform 1 0 31188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1676037725
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1676037725
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_370
timestamp 1676037725
transform 1 0 35144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_378
timestamp 1676037725
transform 1 0 35880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_382
timestamp 1676037725
transform 1 0 36248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1676037725
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_399
timestamp 1676037725
transform 1 0 37812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_409
timestamp 1676037725
transform 1 0 38732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1676037725
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_64
timestamp 1676037725
transform 1 0 6992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_77
timestamp 1676037725
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_101
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1676037725
transform 1 0 13248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_194
timestamp 1676037725
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1676037725
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1676037725
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1676037725
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1676037725
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_292
timestamp 1676037725
transform 1 0 27968 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_298
timestamp 1676037725
transform 1 0 28520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_320
timestamp 1676037725
transform 1 0 30544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1676037725
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_346
timestamp 1676037725
transform 1 0 32936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_354
timestamp 1676037725
transform 1 0 33672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_363
timestamp 1676037725
transform 1 0 34500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_367
timestamp 1676037725
transform 1 0 34868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1676037725
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_398
timestamp 1676037725
transform 1 0 37720 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_404
timestamp 1676037725
transform 1 0 38272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_409
timestamp 1676037725
transform 1 0 38732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_11
timestamp 1676037725
transform 1 0 2116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_40
timestamp 1676037725
transform 1 0 4784 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_46
timestamp 1676037725
transform 1 0 5336 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1676037725
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_69
timestamp 1676037725
transform 1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_105
timestamp 1676037725
transform 1 0 10764 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1676037725
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1676037725
transform 1 0 14536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_170
timestamp 1676037725
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_227
timestamp 1676037725
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1676037725
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_288
timestamp 1676037725
transform 1 0 27600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_316
timestamp 1676037725
transform 1 0 30176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_340
timestamp 1676037725
transform 1 0 32384 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_355
timestamp 1676037725
transform 1 0 33764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1676037725
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_388
timestamp 1676037725
transform 1 0 36800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_395
timestamp 1676037725
transform 1 0 37444 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_403
timestamp 1676037725
transform 1 0 38180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_409
timestamp 1676037725
transform 1 0 38732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_9
timestamp 1676037725
transform 1 0 1932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_17
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_67
timestamp 1676037725
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_80
timestamp 1676037725
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1676037725
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1676037725
transform 1 0 11960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1676037725
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1676037725
transform 1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_203
timestamp 1676037725
transform 1 0 19780 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1676037725
transform 1 0 20516 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1676037725
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1676037725
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_250
timestamp 1676037725
transform 1 0 24104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_263
timestamp 1676037725
transform 1 0 25300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1676037725
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_288
timestamp 1676037725
transform 1 0 27600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_301
timestamp 1676037725
transform 1 0 28796 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_307
timestamp 1676037725
transform 1 0 29348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1676037725
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_360
timestamp 1676037725
transform 1 0 34224 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_377
timestamp 1676037725
transform 1 0 35788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp 1676037725
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_398
timestamp 1676037725
transform 1 0 37720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1676037725
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_38
timestamp 1676037725
transform 1 0 4600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1676037725
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_75
timestamp 1676037725
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1676037725
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_108
timestamp 1676037725
transform 1 0 11040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1676037725
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_150
timestamp 1676037725
transform 1 0 14904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_175
timestamp 1676037725
transform 1 0 17204 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_183
timestamp 1676037725
transform 1 0 17940 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1676037725
transform 1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1676037725
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1676037725
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_264
timestamp 1676037725
transform 1 0 25392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_290
timestamp 1676037725
transform 1 0 27784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1676037725
transform 1 0 31556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1676037725
transform 1 0 31924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp 1676037725
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_371
timestamp 1676037725
transform 1 0 35236 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_381
timestamp 1676037725
transform 1 0 36156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_388
timestamp 1676037725
transform 1 0 36800 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1676037725
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_402
timestamp 1676037725
transform 1 0 38088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_409
timestamp 1676037725
transform 1 0 38732 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1676037725
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_44
timestamp 1676037725
transform 1 0 5152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_79
timestamp 1676037725
transform 1 0 8372 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1676037725
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1676037725
transform 1 0 10028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1676037725
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_142
timestamp 1676037725
transform 1 0 14168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1676037725
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1676037725
transform 1 0 20884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_238
timestamp 1676037725
transform 1 0 23000 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_251
timestamp 1676037725
transform 1 0 24196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_257
timestamp 1676037725
transform 1 0 24748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1676037725
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_290
timestamp 1676037725
transform 1 0 27784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_314
timestamp 1676037725
transform 1 0 29992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_327
timestamp 1676037725
transform 1 0 31188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1676037725
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_343
timestamp 1676037725
transform 1 0 32660 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_347
timestamp 1676037725
transform 1 0 33028 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_368
timestamp 1676037725
transform 1 0 34960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_381
timestamp 1676037725
transform 1 0 36156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1676037725
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_398
timestamp 1676037725
transform 1 0 37720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1676037725
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1676037725
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1676037725
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_108
timestamp 1676037725
transform 1 0 11040 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_116
timestamp 1676037725
transform 1 0 11776 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1676037725
transform 1 0 15272 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_178
timestamp 1676037725
transform 1 0 17480 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_184
timestamp 1676037725
transform 1 0 18032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_204
timestamp 1676037725
transform 1 0 19872 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_217
timestamp 1676037725
transform 1 0 21068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_241
timestamp 1676037725
transform 1 0 23276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1676037725
transform 1 0 25944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1676037725
transform 1 0 26312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_285
timestamp 1676037725
transform 1 0 27324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_298
timestamp 1676037725
transform 1 0 28520 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1676037725
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_320
timestamp 1676037725
transform 1 0 30544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_341
timestamp 1676037725
transform 1 0 32476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1676037725
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_372
timestamp 1676037725
transform 1 0 35328 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_408
timestamp 1676037725
transform 1 0 38640 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_22
timestamp 1676037725
transform 1 0 3128 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1676037725
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp 1676037725
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 1676037725
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_129
timestamp 1676037725
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1676037725
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_182
timestamp 1676037725
transform 1 0 17848 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_206
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1676037725
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_236
timestamp 1676037725
transform 1 0 22816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1676037725
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_257
timestamp 1676037725
transform 1 0 24748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1676037725
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_303
timestamp 1676037725
transform 1 0 28980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_309
timestamp 1676037725
transform 1 0 29532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_330
timestamp 1676037725
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_348
timestamp 1676037725
transform 1 0 33120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_352
timestamp 1676037725
transform 1 0 33488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_360
timestamp 1676037725
transform 1 0 34224 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_384
timestamp 1676037725
transform 1 0 36432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_404
timestamp 1676037725
transform 1 0 38272 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_410
timestamp 1676037725
transform 1 0 38824 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1676037725
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_13
timestamp 1676037725
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1676037725
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_91
timestamp 1676037725
transform 1 0 9476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_104
timestamp 1676037725
transform 1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1676037725
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 1676037725
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_161
timestamp 1676037725
transform 1 0 15916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_169
timestamp 1676037725
transform 1 0 16652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1676037725
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp 1676037725
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_213
timestamp 1676037725
transform 1 0 20700 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1676037725
transform 1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_284
timestamp 1676037725
transform 1 0 27232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_296
timestamp 1676037725
transform 1 0 28336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1676037725
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_315
timestamp 1676037725
transform 1 0 30084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_328
timestamp 1676037725
transform 1 0 31280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_339
timestamp 1676037725
transform 1 0 32292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_354
timestamp 1676037725
transform 1 0 33672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1676037725
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_376
timestamp 1676037725
transform 1 0 35696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_383
timestamp 1676037725
transform 1 0 36340 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_387
timestamp 1676037725
transform 1 0 36708 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_409
timestamp 1676037725
transform 1 0 38732 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1676037725
transform 1 0 2392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_25
timestamp 1676037725
transform 1 0 3404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1676037725
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1676037725
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_100
timestamp 1676037725
transform 1 0 10304 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_106
timestamp 1676037725
transform 1 0 10856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_124
timestamp 1676037725
transform 1 0 12512 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1676037725
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1676037725
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1676037725
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_194
timestamp 1676037725
transform 1 0 18952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1676037725
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_238
timestamp 1676037725
transform 1 0 23000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_251
timestamp 1676037725
transform 1 0 24196 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_255
timestamp 1676037725
transform 1 0 24564 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1676037725
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_292
timestamp 1676037725
transform 1 0 27968 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_298
timestamp 1676037725
transform 1 0 28520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_320
timestamp 1676037725
transform 1 0 30544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1676037725
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_354
timestamp 1676037725
transform 1 0 33672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_363
timestamp 1676037725
transform 1 0 34500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_369
timestamp 1676037725
transform 1 0 35052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1676037725
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_404
timestamp 1676037725
transform 1 0 38272 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_410
timestamp 1676037725
transform 1 0 38824 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1676037725
transform 1 0 2392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1676037725
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_37
timestamp 1676037725
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_50
timestamp 1676037725
transform 1 0 5704 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1676037725
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_96
timestamp 1676037725
transform 1 0 9936 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1676037725
transform 1 0 10672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1676037725
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1676037725
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_146
timestamp 1676037725
transform 1 0 14536 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1676037725
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_174
timestamp 1676037725
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_183
timestamp 1676037725
transform 1 0 17940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_236
timestamp 1676037725
transform 1 0 22816 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 1676037725
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_264
timestamp 1676037725
transform 1 0 25392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_275
timestamp 1676037725
transform 1 0 26404 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_302
timestamp 1676037725
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_331
timestamp 1676037725
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_355
timestamp 1676037725
transform 1 0 33764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1676037725
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_375
timestamp 1676037725
transform 1 0 35604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_400
timestamp 1676037725
transform 1 0 37904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_404
timestamp 1676037725
transform 1 0 38272 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_409
timestamp 1676037725
transform 1 0 38732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_28
timestamp 1676037725
transform 1 0 3680 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_68
timestamp 1676037725
transform 1 0 7360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1676037725
transform 1 0 8096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_101
timestamp 1676037725
transform 1 0 10396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_132
timestamp 1676037725
transform 1 0 13248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_140
timestamp 1676037725
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_150
timestamp 1676037725
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_194
timestamp 1676037725
transform 1 0 18952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_207
timestamp 1676037725
transform 1 0 20148 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_236
timestamp 1676037725
transform 1 0 22816 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_246
timestamp 1676037725
transform 1 0 23736 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_254
timestamp 1676037725
transform 1 0 24472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1676037725
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_304
timestamp 1676037725
transform 1 0 29072 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1676037725
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_348
timestamp 1676037725
transform 1 0 33120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_365
timestamp 1676037725
transform 1 0 34684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_375
timestamp 1676037725
transform 1 0 35604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1676037725
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_404
timestamp 1676037725
transform 1 0 38272 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_410
timestamp 1676037725
transform 1 0 38824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1676037725
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_52
timestamp 1676037725
transform 1 0 5888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_58
timestamp 1676037725
transform 1 0 6440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_68
timestamp 1676037725
transform 1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1676037725
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1676037725
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1676037725
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_123
timestamp 1676037725
transform 1 0 12420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1676037725
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_179
timestamp 1676037725
transform 1 0 17572 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_207
timestamp 1676037725
transform 1 0 20148 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1676037725
transform 1 0 22356 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_275
timestamp 1676037725
transform 1 0 26404 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_283
timestamp 1676037725
transform 1 0 27140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1676037725
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_318
timestamp 1676037725
transform 1 0 30360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_342
timestamp 1676037725
transform 1 0 32568 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_350
timestamp 1676037725
transform 1 0 33304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1676037725
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_376
timestamp 1676037725
transform 1 0 35696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_383
timestamp 1676037725
transform 1 0 36340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_387
timestamp 1676037725
transform 1 0 36708 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_409
timestamp 1676037725
transform 1 0 38732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_9
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_13
timestamp 1676037725
transform 1 0 2300 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_34
timestamp 1676037725
transform 1 0 4232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1676037725
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 1676037725
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_119
timestamp 1676037725
transform 1 0 12052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1676037725
transform 1 0 13248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_158
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_162
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_184
timestamp 1676037725
transform 1 0 18032 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_190
timestamp 1676037725
transform 1 0 18584 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_211
timestamp 1676037725
transform 1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_245
timestamp 1676037725
transform 1 0 23644 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_266
timestamp 1676037725
transform 1 0 25576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_270
timestamp 1676037725
transform 1 0 25944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_296
timestamp 1676037725
transform 1 0 28336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_310
timestamp 1676037725
transform 1 0 29624 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1676037725
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_345
timestamp 1676037725
transform 1 0 32844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_370
timestamp 1676037725
transform 1 0 35144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_383
timestamp 1676037725
transform 1 0 36340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_398
timestamp 1676037725
transform 1 0 37720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_9
timestamp 1676037725
transform 1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1676037725
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_21
timestamp 1676037725
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_42
timestamp 1676037725
transform 1 0 4968 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_51
timestamp 1676037725
transform 1 0 5796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1676037725
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1676037725
transform 1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_113
timestamp 1676037725
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_117
timestamp 1676037725
transform 1 0 11868 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1676037725
transform 1 0 12604 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_146
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_150
timestamp 1676037725
transform 1 0 14904 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_160
timestamp 1676037725
transform 1 0 15824 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1676037725
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_208
timestamp 1676037725
transform 1 0 20240 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_235
timestamp 1676037725
transform 1 0 22724 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1676037725
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_260
timestamp 1676037725
transform 1 0 25024 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_276
timestamp 1676037725
transform 1 0 26496 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_297
timestamp 1676037725
transform 1 0 28428 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1676037725
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1676037725
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_327
timestamp 1676037725
transform 1 0 31188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_336
timestamp 1676037725
transform 1 0 32016 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_347
timestamp 1676037725
transform 1 0 33028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_358
timestamp 1676037725
transform 1 0 34040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_390
timestamp 1676037725
transform 1 0 36984 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_397
timestamp 1676037725
transform 1 0 37628 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_409
timestamp 1676037725
transform 1 0 38732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_13
timestamp 1676037725
transform 1 0 2300 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 1676037725
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_67
timestamp 1676037725
transform 1 0 7268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_94
timestamp 1676037725
transform 1 0 9752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_121
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_147
timestamp 1676037725
transform 1 0 14628 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1676037725
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_180
timestamp 1676037725
transform 1 0 17664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_204
timestamp 1676037725
transform 1 0 19872 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1676037725
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_257
timestamp 1676037725
transform 1 0 24748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_266
timestamp 1676037725
transform 1 0 25576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1676037725
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_292
timestamp 1676037725
transform 1 0 27968 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_300
timestamp 1676037725
transform 1 0 28704 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_321
timestamp 1676037725
transform 1 0 30636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1676037725
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_359
timestamp 1676037725
transform 1 0 34132 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_383
timestamp 1676037725
transform 1 0 36340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1676037725
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_398
timestamp 1676037725
transform 1 0 37720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_11
timestamp 1676037725
transform 1 0 2116 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_51
timestamp 1676037725
transform 1 0 5796 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_55
timestamp 1676037725
transform 1 0 6164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1676037725
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1676037725
transform 1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_75
timestamp 1676037725
transform 1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_107
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_125
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_164
timestamp 1676037725
transform 1 0 16192 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_179
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1676037725
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_206
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_216
timestamp 1676037725
transform 1 0 20976 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_241
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_270
timestamp 1676037725
transform 1 0 25944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_281
timestamp 1676037725
transform 1 0 26956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_295
timestamp 1676037725
transform 1 0 28244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_302
timestamp 1676037725
transform 1 0 28888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_314
timestamp 1676037725
transform 1 0 29992 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_331
timestamp 1676037725
transform 1 0 31556 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_338
timestamp 1676037725
transform 1 0 32200 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_370
timestamp 1676037725
transform 1 0 35144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_384
timestamp 1676037725
transform 1 0 36432 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_391
timestamp 1676037725
transform 1 0 37076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_395
timestamp 1676037725
transform 1 0 37444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1676037725
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_409
timestamp 1676037725
transform 1 0 38732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_10
timestamp 1676037725
transform 1 0 2024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_35
timestamp 1676037725
transform 1 0 4324 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_43
timestamp 1676037725
transform 1 0 5060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_68
timestamp 1676037725
transform 1 0 7360 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_74
timestamp 1676037725
transform 1 0 7912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1676037725
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_89
timestamp 1676037725
transform 1 0 9292 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_102
timestamp 1676037725
transform 1 0 10488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_106
timestamp 1676037725
transform 1 0 10856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_124
timestamp 1676037725
transform 1 0 12512 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1676037725
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_182
timestamp 1676037725
transform 1 0 17848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1676037725
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_202
timestamp 1676037725
transform 1 0 19688 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_215
timestamp 1676037725
transform 1 0 20884 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_234
timestamp 1676037725
transform 1 0 22632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_238
timestamp 1676037725
transform 1 0 23000 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_259
timestamp 1676037725
transform 1 0 24932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_272
timestamp 1676037725
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_303
timestamp 1676037725
transform 1 0 28980 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_307
timestamp 1676037725
transform 1 0 29348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_313
timestamp 1676037725
transform 1 0 29900 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_328
timestamp 1676037725
transform 1 0 31280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_352
timestamp 1676037725
transform 1 0 33488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_359
timestamp 1676037725
transform 1 0 34132 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_387
timestamp 1676037725
transform 1 0 36708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_404
timestamp 1676037725
transform 1 0 38272 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_410
timestamp 1676037725
transform 1 0 38824 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_12
timestamp 1676037725
transform 1 0 2208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_19
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1676037725
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_51
timestamp 1676037725
transform 1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_55
timestamp 1676037725
transform 1 0 6164 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_59
timestamp 1676037725
transform 1 0 6532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_72
timestamp 1676037725
transform 1 0 7728 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_78
timestamp 1676037725
transform 1 0 8280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_96
timestamp 1676037725
transform 1 0 9936 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_103
timestamp 1676037725
transform 1 0 10580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1676037725
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1676037725
transform 1 0 12788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_146
timestamp 1676037725
transform 1 0 14536 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1676037725
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_161
timestamp 1676037725
transform 1 0 15916 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_171
timestamp 1676037725
transform 1 0 16836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_182
timestamp 1676037725
transform 1 0 17848 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1676037725
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1676037725
transform 1 0 20884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_228
timestamp 1676037725
transform 1 0 22080 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_238
timestamp 1676037725
transform 1 0 23000 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_246
timestamp 1676037725
transform 1 0 23736 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1676037725
transform 1 0 24748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_261
timestamp 1676037725
transform 1 0 25116 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_287
timestamp 1676037725
transform 1 0 27508 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 1676037725
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_315
timestamp 1676037725
transform 1 0 30084 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_336
timestamp 1676037725
transform 1 0 32016 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_358
timestamp 1676037725
transform 1 0 34040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_373
timestamp 1676037725
transform 1 0 35420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_383
timestamp 1676037725
transform 1 0 36340 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_390
timestamp 1676037725
transform 1 0 36984 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_398
timestamp 1676037725
transform 1 0 37720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1676037725
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_409
timestamp 1676037725
transform 1 0 38732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_8
timestamp 1676037725
transform 1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_35
timestamp 1676037725
transform 1 0 4324 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_43
timestamp 1676037725
transform 1 0 5060 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_47
timestamp 1676037725
transform 1 0 5428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1676037725
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1676037725
transform 1 0 7176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1676037725
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_89
timestamp 1676037725
transform 1 0 9292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1676037725
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_103
timestamp 1676037725
transform 1 0 10580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_124
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_130
timestamp 1676037725
transform 1 0 13064 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_136
timestamp 1676037725
transform 1 0 13616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_143
timestamp 1676037725
transform 1 0 14260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_157
timestamp 1676037725
transform 1 0 15548 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1676037725
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_233
timestamp 1676037725
transform 1 0 22540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_257
timestamp 1676037725
transform 1 0 24748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_264
timestamp 1676037725
transform 1 0 25392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_268
timestamp 1676037725
transform 1 0 25760 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1676037725
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1676037725
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_299
timestamp 1676037725
transform 1 0 28612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_307
timestamp 1676037725
transform 1 0 29348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1676037725
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_343
timestamp 1676037725
transform 1 0 32660 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_351
timestamp 1676037725
transform 1 0 33396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_358
timestamp 1676037725
transform 1 0 34040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_371
timestamp 1676037725
transform 1 0 35236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1676037725
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_399
timestamp 1676037725
transform 1 0 37812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_406
timestamp 1676037725
transform 1 0 38456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_410
timestamp 1676037725
transform 1 0 38824 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_9
timestamp 1676037725
transform 1 0 1932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_19
timestamp 1676037725
transform 1 0 2852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1676037725
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_47
timestamp 1676037725
transform 1 0 5428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_51
timestamp 1676037725
transform 1 0 5796 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_72
timestamp 1676037725
transform 1 0 7728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_96
timestamp 1676037725
transform 1 0 9936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_103
timestamp 1676037725
transform 1 0 10580 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1676037725
transform 1 0 12604 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1676037725
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_147
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 1676037725
transform 1 0 15548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_171
timestamp 1676037725
transform 1 0 16836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1676037725
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1676037725
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_233
timestamp 1676037725
transform 1 0 22540 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_242
timestamp 1676037725
transform 1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_268
timestamp 1676037725
transform 1 0 25760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_281
timestamp 1676037725
transform 1 0 26956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_294
timestamp 1676037725
transform 1 0 28152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1676037725
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_314
timestamp 1676037725
transform 1 0 29992 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_340
timestamp 1676037725
transform 1 0 32384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_353
timestamp 1676037725
transform 1 0 33580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1676037725
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_387
timestamp 1676037725
transform 1 0 36708 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_395
timestamp 1676037725
transform 1 0 37444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_399
timestamp 1676037725
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_409
timestamp 1676037725
transform 1 0 38732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_28
timestamp 1676037725
transform 1 0 3680 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1676037725
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_74
timestamp 1676037725
transform 1 0 7912 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 1676037725
transform 1 0 9108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1676037725
transform 1 0 10028 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1676037725
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_117
timestamp 1676037725
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_121
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1676037725
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1676037725
transform 1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_180
timestamp 1676037725
transform 1 0 17664 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_188
timestamp 1676037725
transform 1 0 18400 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_249
timestamp 1676037725
transform 1 0 24012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_257
timestamp 1676037725
transform 1 0 24748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_286
timestamp 1676037725
transform 1 0 27416 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_314
timestamp 1676037725
transform 1 0 29992 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_323
timestamp 1676037725
transform 1 0 30820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_327
timestamp 1676037725
transform 1 0 31188 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1676037725
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_348
timestamp 1676037725
transform 1 0 33120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_352
timestamp 1676037725
transform 1 0 33488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_360
timestamp 1676037725
transform 1 0 34224 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_367
timestamp 1676037725
transform 1 0 34868 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_382
timestamp 1676037725
transform 1 0 36248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_386
timestamp 1676037725
transform 1 0 36616 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1676037725
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_398
timestamp 1676037725
transform 1 0 37720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_13
timestamp 1676037725
transform 1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_36
timestamp 1676037725
transform 1 0 4416 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_62
timestamp 1676037725
transform 1 0 6808 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_96
timestamp 1676037725
transform 1 0 9936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_124
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 1676037725
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1676037725
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_184
timestamp 1676037725
transform 1 0 18032 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_234 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22632 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1676037725
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_281
timestamp 1676037725
transform 1 0 26956 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_293
timestamp 1676037725
transform 1 0 28060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_320
timestamp 1676037725
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_324
timestamp 1676037725
transform 1 0 30912 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_346
timestamp 1676037725
transform 1 0 32936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_359
timestamp 1676037725
transform 1 0 34132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_388
timestamp 1676037725
transform 1 0 36800 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_396
timestamp 1676037725
transform 1 0 37536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_403
timestamp 1676037725
transform 1 0 38180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1676037725
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_19
timestamp 1676037725
transform 1 0 2852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_40
timestamp 1676037725
transform 1 0 4784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1676037725
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_66
timestamp 1676037725
transform 1 0 7176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1676037725
transform 1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_80
timestamp 1676037725
transform 1 0 8464 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_101
timestamp 1676037725
transform 1 0 10396 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_124
timestamp 1676037725
transform 1 0 12512 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_132
timestamp 1676037725
transform 1 0 13248 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_144
timestamp 1676037725
transform 1 0 14352 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_233
timestamp 1676037725
transform 1 0 22540 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_262
timestamp 1676037725
transform 1 0 25208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1676037725
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_303
timestamp 1676037725
transform 1 0 28980 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_319
timestamp 1676037725
transform 1 0 30452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_328
timestamp 1676037725
transform 1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_359
timestamp 1676037725
transform 1 0 34132 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1676037725
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_397
timestamp 1676037725
transform 1 0 37628 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_401
timestamp 1676037725
transform 1 0 37996 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_409
timestamp 1676037725
transform 1 0 38732 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_11
timestamp 1676037725
transform 1 0 2116 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1676037725
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_51
timestamp 1676037725
transform 1 0 5796 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_58
timestamp 1676037725
transform 1 0 6440 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_73
timestamp 1676037725
transform 1 0 7820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1676037725
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_90
timestamp 1676037725
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_154
timestamp 1676037725
transform 1 0 15272 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_160
timestamp 1676037725
transform 1 0 15824 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1676037725
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_205
timestamp 1676037725
transform 1 0 19964 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_237
timestamp 1676037725
transform 1 0 22908 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_259
timestamp 1676037725
transform 1 0 24932 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_270
timestamp 1676037725
transform 1 0 25944 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1676037725
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_289
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_295
timestamp 1676037725
transform 1 0 28244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_323
timestamp 1676037725
transform 1 0 30820 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_336
timestamp 1676037725
transform 1 0 32016 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_340
timestamp 1676037725
transform 1 0 32384 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_350
timestamp 1676037725
transform 1 0 33304 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_359
timestamp 1676037725
transform 1 0 34132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_392
timestamp 1676037725
transform 1 0 37168 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_405
timestamp 1676037725
transform 1 0 38364 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_8
timestamp 1676037725
transform 1 0 1840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_32
timestamp 1676037725
transform 1 0 4048 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1676037725
transform 1 0 4784 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_90
timestamp 1676037725
transform 1 0 9384 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_102
timestamp 1676037725
transform 1 0 10488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_106
timestamp 1676037725
transform 1 0 10856 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_128
timestamp 1676037725
transform 1 0 12880 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1676037725
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_177
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_189
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_201
timestamp 1676037725
transform 1 0 19596 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_213
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1676037725
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_259
timestamp 1676037725
transform 1 0 24932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_271
timestamp 1676037725
transform 1 0 26036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_285
timestamp 1676037725
transform 1 0 27324 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_306
timestamp 1676037725
transform 1 0 29256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1676037725
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_344
timestamp 1676037725
transform 1 0 32752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_369
timestamp 1676037725
transform 1 0 35052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_382
timestamp 1676037725
transform 1 0 36248 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1676037725
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_398
timestamp 1676037725
transform 1 0 37720 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_410
timestamp 1676037725
transform 1 0 38824 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_19
timestamp 1676037725
transform 1 0 2852 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_44
timestamp 1676037725
transform 1 0 5152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1676037725
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_58
timestamp 1676037725
transform 1 0 6440 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_70
timestamp 1676037725
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_130
timestamp 1676037725
transform 1 0 13064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_134
timestamp 1676037725
transform 1 0 13432 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_178
timestamp 1676037725
transform 1 0 17480 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185
timestamp 1676037725
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1676037725
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_215
timestamp 1676037725
transform 1 0 20884 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1676037725
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1676037725
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_266
timestamp 1676037725
transform 1 0 25576 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_274
timestamp 1676037725
transform 1 0 26312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_281
timestamp 1676037725
transform 1 0 26956 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1676037725
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_315
timestamp 1676037725
transform 1 0 30084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_325
timestamp 1676037725
transform 1 0 31004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_340
timestamp 1676037725
transform 1 0 32384 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_353
timestamp 1676037725
transform 1 0 33580 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_374
timestamp 1676037725
transform 1 0 35512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_381
timestamp 1676037725
transform 1 0 36156 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_388
timestamp 1676037725
transform 1 0 36800 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_400
timestamp 1676037725
transform 1 0 37904 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_408
timestamp 1676037725
transform 1 0 38640 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_8
timestamp 1676037725
transform 1 0 1840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_36
timestamp 1676037725
transform 1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1676037725
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_80
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_92
timestamp 1676037725
transform 1 0 9568 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_104
timestamp 1676037725
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1676037725
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_194
timestamp 1676037725
transform 1 0 18952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_243
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_250
timestamp 1676037725
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_265
timestamp 1676037725
transform 1 0 25484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1676037725
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_287
timestamp 1676037725
transform 1 0 27508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_299
timestamp 1676037725
transform 1 0 28612 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_307
timestamp 1676037725
transform 1 0 29348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_319
timestamp 1676037725
transform 1 0 30452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_347
timestamp 1676037725
transform 1 0 33028 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_364
timestamp 1676037725
transform 1 0 34592 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_377
timestamp 1676037725
transform 1 0 35788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1676037725
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_409
timestamp 1676037725
transform 1 0 38732 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1676037725
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_13
timestamp 1676037725
transform 1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1676037725
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_157
timestamp 1676037725
transform 1 0 15548 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_178
timestamp 1676037725
transform 1 0 17480 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1676037725
transform 1 0 19964 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_213
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_226
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_273
timestamp 1676037725
transform 1 0 26220 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_287
timestamp 1676037725
transform 1 0 27508 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_299
timestamp 1676037725
transform 1 0 28612 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1676037725
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_314
timestamp 1676037725
transform 1 0 29992 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_322
timestamp 1676037725
transform 1 0 30728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_348
timestamp 1676037725
transform 1 0 33120 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_354
timestamp 1676037725
transform 1 0 33672 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1676037725
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1676037725
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_401
timestamp 1676037725
transform 1 0 37996 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_409
timestamp 1676037725
transform 1 0 38732 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_38
timestamp 1676037725
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1676037725
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_175
timestamp 1676037725
transform 1 0 17204 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_183
timestamp 1676037725
transform 1 0 17940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_195
timestamp 1676037725
transform 1 0 19044 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1676037725
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1676037725
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1676037725
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_251
timestamp 1676037725
transform 1 0 24196 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_289
timestamp 1676037725
transform 1 0 27692 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_301
timestamp 1676037725
transform 1 0 28796 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_321
timestamp 1676037725
transform 1 0 30636 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1676037725
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1676037725
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 1676037725
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_398
timestamp 1676037725
transform 1 0 37720 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_410
timestamp 1676037725
transform 1 0 38824 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_9
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_52
timestamp 1676037725
transform 1 0 5888 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_71
timestamp 1676037725
transform 1 0 7636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_117
timestamp 1676037725
transform 1 0 11868 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_122
timestamp 1676037725
transform 1 0 12328 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1676037725
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1676037725
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_203
timestamp 1676037725
transform 1 0 19780 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1676037725
transform 1 0 20424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_234
timestamp 1676037725
transform 1 0 22632 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1676037725
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1676037725
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_257
timestamp 1676037725
transform 1 0 24748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_267
timestamp 1676037725
transform 1 0 25668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_277
timestamp 1676037725
transform 1 0 26588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_290
timestamp 1676037725
transform 1 0 27784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_297
timestamp 1676037725
transform 1 0 28428 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_305
timestamp 1676037725
transform 1 0 29164 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_317
timestamp 1676037725
transform 1 0 30268 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_329
timestamp 1676037725
transform 1 0 31372 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_337
timestamp 1676037725
transform 1 0 32108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1676037725
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_373
timestamp 1676037725
transform 1 0 35420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_387
timestamp 1676037725
transform 1 0 36708 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_400
timestamp 1676037725
transform 1 0 37904 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_408
timestamp 1676037725
transform 1 0 38640 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_38
timestamp 1676037725
transform 1 0 4600 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_46
timestamp 1676037725
transform 1 0 5336 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_119
timestamp 1676037725
transform 1 0 12052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_144
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_155
timestamp 1676037725
transform 1 0 15364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_177
timestamp 1676037725
transform 1 0 17388 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_201
timestamp 1676037725
transform 1 0 19596 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_209
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_251
timestamp 1676037725
transform 1 0 24196 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1676037725
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1676037725
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_317
timestamp 1676037725
transform 1 0 30268 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_321
timestamp 1676037725
transform 1 0 30636 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1676037725
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1676037725
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_376
timestamp 1676037725
transform 1 0 35696 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1676037725
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1676037725
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_45
timestamp 1676037725
transform 1 0 5244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_48
timestamp 1676037725
transform 1 0 5520 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_56
timestamp 1676037725
transform 1 0 6256 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_68
timestamp 1676037725
transform 1 0 7360 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1676037725
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_149
timestamp 1676037725
transform 1 0 14812 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_161
timestamp 1676037725
transform 1 0 15916 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_173
timestamp 1676037725
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_185
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_205
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1676037725
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1676037725
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_238
timestamp 1676037725
transform 1 0 23000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1676037725
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1676037725
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1676037725
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_321
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_327
timestamp 1676037725
transform 1 0 31188 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_348
timestamp 1676037725
transform 1 0 33120 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1676037725
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_401
timestamp 1676037725
transform 1 0 37996 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_409
timestamp 1676037725
transform 1 0 38732 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_11
timestamp 1676037725
transform 1 0 2116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_33
timestamp 1676037725
transform 1 0 4140 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_40
timestamp 1676037725
transform 1 0 4784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1676037725
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_123
timestamp 1676037725
transform 1 0 12420 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_135
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_147
timestamp 1676037725
transform 1 0 14628 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1676037725
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_231
timestamp 1676037725
transform 1 0 22356 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_238
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_244
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_248
timestamp 1676037725
transform 1 0 23920 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_260
timestamp 1676037725
transform 1 0 25024 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1676037725
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_292
timestamp 1676037725
transform 1 0 27968 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_309
timestamp 1676037725
transform 1 0 29532 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_321
timestamp 1676037725
transform 1 0 30636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1676037725
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_345
timestamp 1676037725
transform 1 0 32844 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_357
timestamp 1676037725
transform 1 0 33948 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_369
timestamp 1676037725
transform 1 0 35052 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_377
timestamp 1676037725
transform 1 0 35788 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_383
timestamp 1676037725
transform 1 0 36340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1676037725
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_11
timestamp 1676037725
transform 1 0 2116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 1676037725
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_34
timestamp 1676037725
transform 1 0 4232 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_46
timestamp 1676037725
transform 1 0 5336 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_58
timestamp 1676037725
transform 1 0 6440 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_70
timestamp 1676037725
transform 1 0 7544 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_112
timestamp 1676037725
transform 1 0 11408 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_120
timestamp 1676037725
transform 1 0 12144 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_281
timestamp 1676037725
transform 1 0 26956 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_289
timestamp 1676037725
transform 1 0 27692 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_299
timestamp 1676037725
transform 1 0 28612 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_316
timestamp 1676037725
transform 1 0 30176 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_324
timestamp 1676037725
transform 1 0 30912 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_328
timestamp 1676037725
transform 1 0 31280 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_340
timestamp 1676037725
transform 1 0 32384 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_352
timestamp 1676037725
transform 1 0 33488 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_390
timestamp 1676037725
transform 1 0 36984 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_402
timestamp 1676037725
transform 1 0 38088 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_409
timestamp 1676037725
transform 1 0 38732 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_36
timestamp 1676037725
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1676037725
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_132
timestamp 1676037725
transform 1 0 13248 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_144
timestamp 1676037725
transform 1 0 14352 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_156
timestamp 1676037725
transform 1 0 15456 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_192
timestamp 1676037725
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_204
timestamp 1676037725
transform 1 0 19872 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1676037725
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1676037725
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_249
timestamp 1676037725
transform 1 0 24012 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_315
timestamp 1676037725
transform 1 0 30084 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1676037725
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1676037725
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_373
timestamp 1676037725
transform 1 0 35420 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_379
timestamp 1676037725
transform 1 0 35972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_405
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_40
timestamp 1676037725
transform 1 0 4784 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_52
timestamp 1676037725
transform 1 0 5888 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_64
timestamp 1676037725
transform 1 0 6992 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_76
timestamp 1676037725
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_103
timestamp 1676037725
transform 1 0 10580 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_124
timestamp 1676037725
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1676037725
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_152
timestamp 1676037725
transform 1 0 15088 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_170
timestamp 1676037725
transform 1 0 16744 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_182
timestamp 1676037725
transform 1 0 17848 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1676037725
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1676037725
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_289
timestamp 1676037725
transform 1 0 27692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_297
timestamp 1676037725
transform 1 0 28428 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1676037725
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1676037725
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_315
timestamp 1676037725
transform 1 0 30084 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_319
timestamp 1676037725
transform 1 0 30452 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_336
timestamp 1676037725
transform 1 0 32016 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_349
timestamp 1676037725
transform 1 0 33212 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1676037725
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_409
timestamp 1676037725
transform 1 0 38732 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_9
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_13
timestamp 1676037725
transform 1 0 2300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_25
timestamp 1676037725
transform 1 0 3404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_30
timestamp 1676037725
transform 1 0 3864 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_36
timestamp 1676037725
transform 1 0 4416 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_42
timestamp 1676037725
transform 1 0 4968 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_48
timestamp 1676037725
transform 1 0 5520 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_97
timestamp 1676037725
transform 1 0 10028 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_134
timestamp 1676037725
transform 1 0 13432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_138
timestamp 1676037725
transform 1 0 13800 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1676037725
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_181
timestamp 1676037725
transform 1 0 17756 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_196
timestamp 1676037725
transform 1 0 19136 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1676037725
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_245
timestamp 1676037725
transform 1 0 23644 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_257
timestamp 1676037725
transform 1 0 24748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1676037725
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1676037725
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1676037725
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_350
timestamp 1676037725
transform 1 0 33304 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_362
timestamp 1676037725
transform 1 0 34408 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_374
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_386
timestamp 1676037725
transform 1 0 36616 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_11
timestamp 1676037725
transform 1 0 2116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1676037725
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_66
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_78
timestamp 1676037725
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_92
timestamp 1676037725
transform 1 0 9568 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_100
timestamp 1676037725
transform 1 0 10304 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_112
timestamp 1676037725
transform 1 0 11408 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_124
timestamp 1676037725
transform 1 0 12512 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_128
timestamp 1676037725
transform 1 0 12880 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_146
timestamp 1676037725
transform 1 0 14536 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_158
timestamp 1676037725
transform 1 0 15640 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_182
timestamp 1676037725
transform 1 0 17848 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_268
timestamp 1676037725
transform 1 0 25760 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_280
timestamp 1676037725
transform 1 0 26864 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_292
timestamp 1676037725
transform 1 0 27968 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1676037725
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_321
timestamp 1676037725
transform 1 0 30636 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_329
timestamp 1676037725
transform 1 0 31372 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_337
timestamp 1676037725
transform 1 0 32108 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_349
timestamp 1676037725
transform 1 0 33212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_401
timestamp 1676037725
transform 1 0 37996 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_409
timestamp 1676037725
transform 1 0 38732 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_45
timestamp 1676037725
transform 1 0 5244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1676037725
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_68
timestamp 1676037725
transform 1 0 7360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_72
timestamp 1676037725
transform 1 0 7728 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_82
timestamp 1676037725
transform 1 0 8648 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_95
timestamp 1676037725
transform 1 0 9844 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_107
timestamp 1676037725
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_132
timestamp 1676037725
transform 1 0 13248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1676037725
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_155
timestamp 1676037725
transform 1 0 15364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_187
timestamp 1676037725
transform 1 0 18308 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_199
timestamp 1676037725
transform 1 0 19412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_211
timestamp 1676037725
transform 1 0 20516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_249
timestamp 1676037725
transform 1 0 24012 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_257
timestamp 1676037725
transform 1 0 24748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1676037725
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1676037725
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1676037725
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_348
timestamp 1676037725
transform 1 0 33120 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_360
timestamp 1676037725
transform 1 0 34224 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_376
timestamp 1676037725
transform 1 0 35696 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1676037725
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_14
timestamp 1676037725
transform 1 0 2392 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_49
timestamp 1676037725
transform 1 0 5612 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_72
timestamp 1676037725
transform 1 0 7728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_76
timestamp 1676037725
transform 1 0 8096 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1676037725
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_94
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_106
timestamp 1676037725
transform 1 0 10856 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_124
timestamp 1676037725
transform 1 0 12512 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1676037725
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_152
timestamp 1676037725
transform 1 0 15088 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_181
timestamp 1676037725
transform 1 0 17756 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1676037725
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1676037725
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1676037725
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_273
timestamp 1676037725
transform 1 0 26220 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_288
timestamp 1676037725
transform 1 0 27600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_292
timestamp 1676037725
transform 1 0 27968 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_296
timestamp 1676037725
transform 1 0 28336 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_333
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_350
timestamp 1676037725
transform 1 0 33304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_379
timestamp 1676037725
transform 1 0 35972 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_392
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_404
timestamp 1676037725
transform 1 0 38272 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_410
timestamp 1676037725
transform 1 0 38824 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_134
timestamp 1676037725
transform 1 0 13432 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_143
timestamp 1676037725
transform 1 0 14260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_159
timestamp 1676037725
transform 1 0 15732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_177
timestamp 1676037725
transform 1 0 17388 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_188
timestamp 1676037725
transform 1 0 18400 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_200
timestamp 1676037725
transform 1 0 19504 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_212
timestamp 1676037725
transform 1 0 20608 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_257
timestamp 1676037725
transform 1 0 24748 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_263
timestamp 1676037725
transform 1 0 25300 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_275
timestamp 1676037725
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_305
timestamp 1676037725
transform 1 0 29164 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_313
timestamp 1676037725
transform 1 0 29900 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_319
timestamp 1676037725
transform 1 0 30452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1676037725
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_360
timestamp 1676037725
transform 1 0 34224 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_375
timestamp 1676037725
transform 1 0 35604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1676037725
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_399
timestamp 1676037725
transform 1 0 37812 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_409
timestamp 1676037725
transform 1 0 38732 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_9
timestamp 1676037725
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1676037725
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_61
timestamp 1676037725
transform 1 0 6716 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_71
timestamp 1676037725
transform 1 0 7636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1676037725
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_175
timestamp 1676037725
transform 1 0 17204 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_181
timestamp 1676037725
transform 1 0 17756 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1676037725
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1676037725
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_300
timestamp 1676037725
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1676037725
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_333
timestamp 1676037725
transform 1 0 31740 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_341
timestamp 1676037725
transform 1 0 32476 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_351
timestamp 1676037725
transform 1 0 33396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1676037725
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_377
timestamp 1676037725
transform 1 0 35788 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1676037725
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_401
timestamp 1676037725
transform 1 0 37996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_409
timestamp 1676037725
transform 1 0 38732 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_9
timestamp 1676037725
transform 1 0 1932 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_21
timestamp 1676037725
transform 1 0 3036 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_33
timestamp 1676037725
transform 1 0 4140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_45
timestamp 1676037725
transform 1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1676037725
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_134
timestamp 1676037725
transform 1 0 13432 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_146
timestamp 1676037725
transform 1 0 14536 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1676037725
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_162
timestamp 1676037725
transform 1 0 16008 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1676037725
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_175
timestamp 1676037725
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_188
timestamp 1676037725
transform 1 0 18400 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_200
timestamp 1676037725
transform 1 0 19504 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_212
timestamp 1676037725
transform 1 0 20608 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1676037725
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_309
timestamp 1676037725
transform 1 0 29532 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_321
timestamp 1676037725
transform 1 0 30636 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1676037725
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1676037725
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1676037725
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1676037725
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1676037725
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1676037725
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_399
timestamp 1676037725
transform 1 0 37812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_409
timestamp 1676037725
transform 1 0 38732 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1676037725
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_16
timestamp 1676037725
transform 1 0 2576 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1676037725
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_37
timestamp 1676037725
transform 1 0 4508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_49
timestamp 1676037725
transform 1 0 5612 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_55
timestamp 1676037725
transform 1 0 6164 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_57
timestamp 1676037725
transform 1 0 6348 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_93
timestamp 1676037725
transform 1 0 9660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_105
timestamp 1676037725
transform 1 0 10764 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_111
timestamp 1676037725
transform 1 0 11316 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_113
timestamp 1676037725
transform 1 0 11500 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_119
timestamp 1676037725
transform 1 0 12052 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_127
timestamp 1676037725
transform 1 0 12788 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1676037725
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_149
timestamp 1676037725
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_156
timestamp 1676037725
transform 1 0 15456 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_169
timestamp 1676037725
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_175
timestamp 1676037725
transform 1 0 17204 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_183
timestamp 1676037725
transform 1 0 17940 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_191
timestamp 1676037725
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_205
timestamp 1676037725
transform 1 0 19964 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_210
timestamp 1676037725
transform 1 0 20424 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_222
timestamp 1676037725
transform 1 0 21528 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_225
timestamp 1676037725
transform 1 0 21804 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_231
timestamp 1676037725
transform 1 0 22356 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_239
timestamp 1676037725
transform 1 0 23092 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_247
timestamp 1676037725
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_261
timestamp 1676037725
transform 1 0 25116 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_268
timestamp 1676037725
transform 1 0 25760 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_281
timestamp 1676037725
transform 1 0 26956 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_287
timestamp 1676037725
transform 1 0 27508 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_293
timestamp 1676037725
transform 1 0 28060 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1676037725
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_317
timestamp 1676037725
transform 1 0 30268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_327
timestamp 1676037725
transform 1 0 31188 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_335
timestamp 1676037725
transform 1 0 31924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_337
timestamp 1676037725
transform 1 0 32108 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_343
timestamp 1676037725
transform 1 0 32660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_355
timestamp 1676037725
transform 1 0 33764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1676037725
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_373
timestamp 1676037725
transform 1 0 35420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_387
timestamp 1676037725
transform 1 0 36708 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_391
timestamp 1676037725
transform 1 0 37076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_393
timestamp 1676037725
transform 1 0 37260 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_399
timestamp 1676037725
transform 1 0 37812 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_409
timestamp 1676037725
transform 1 0 38732 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 39192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 39192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 39192 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 39192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 39192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 39192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 39192 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 39192 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 39192 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 39192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 39192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 39192 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 39192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 39192 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 39192 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 39192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 39192 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 39192 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 39192 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 39192 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 39192 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 39192 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 39192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 39192 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 39192 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 39192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 39192 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 39192 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 39192 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 39192 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 39192 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 39192 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 39192 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 39192 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 39192 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 39192 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 39192 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 39192 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 39192 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 39192 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 39192 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 39192 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 39192 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 39192 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 39192 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 11408 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 21712 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 26864 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 32016 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 37168 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _0512_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0513_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13616 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0514_
timestamp 1676037725
transform 1 0 31004 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0515_
timestamp 1676037725
transform 1 0 2668 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0516_
timestamp 1676037725
transform 1 0 19872 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0517_
timestamp 1676037725
transform 1 0 32292 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0518_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0519_
timestamp 1676037725
transform 1 0 25852 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0520_
timestamp 1676037725
transform 1 0 7820 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0521_
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0522_
timestamp 1676037725
transform 1 0 8280 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1676037725
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0524_
timestamp 1676037725
transform 1 0 2668 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0525_
timestamp 1676037725
transform 1 0 7544 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0526_
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0527_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0528_
timestamp 1676037725
transform 1 0 2668 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0529_
timestamp 1676037725
transform 1 0 9844 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0530_
timestamp 1676037725
transform 1 0 4968 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0531_
timestamp 1676037725
transform 1 0 18124 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0532_
timestamp 1676037725
transform 1 0 18124 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0533_
timestamp 1676037725
transform 1 0 33120 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0534_
timestamp 1676037725
transform 1 0 23368 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0535_
timestamp 1676037725
transform 1 0 23092 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0536_
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0537_
timestamp 1676037725
transform 1 0 15548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0538_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0539_
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0540_
timestamp 1676037725
transform 1 0 26956 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0541_
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0542_
timestamp 1676037725
transform 1 0 6348 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0543_
timestamp 1676037725
transform 1 0 30636 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0544_
timestamp 1676037725
transform 1 0 2852 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36340 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0546_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0547_
timestamp 1676037725
transform 1 0 27140 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0548_
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0549_
timestamp 1676037725
transform 1 0 33212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0550_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0551_
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0552_
timestamp 1676037725
transform 1 0 35328 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0553_
timestamp 1676037725
transform 1 0 6808 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0554_
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0555_
timestamp 1676037725
transform 1 0 12144 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0556_
timestamp 1676037725
transform 1 0 32292 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0557_
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 1676037725
transform 1 0 2668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0559_
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0560_
timestamp 1676037725
transform 1 0 29808 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1676037725
transform 1 0 2668 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0562_
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0563_
timestamp 1676037725
transform 1 0 5244 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0564_
timestamp 1676037725
transform 1 0 20700 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0565_
timestamp 1676037725
transform 1 0 17572 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0566_
timestamp 1676037725
transform 1 0 12972 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0567_
timestamp 1676037725
transform 1 0 7360 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0568_
timestamp 1676037725
transform 1 0 28704 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0569_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1676037725
transform 1 0 20240 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0571_
timestamp 1676037725
transform 1 0 10304 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0572_
timestamp 1676037725
transform 1 0 6900 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0573_
timestamp 1676037725
transform 1 0 25668 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0574_
timestamp 1676037725
transform 1 0 29624 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0575_
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0576_
timestamp 1676037725
transform 1 0 32384 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0577_
timestamp 1676037725
transform 1 0 6532 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_4  _0578_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0579_
timestamp 1676037725
transform 1 0 5244 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0580_
timestamp 1676037725
transform 1 0 21252 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0581_
timestamp 1676037725
transform 1 0 28428 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0582_
timestamp 1676037725
transform 1 0 30912 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0583_
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 1676037725
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0585_
timestamp 1676037725
transform 1 0 27140 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0586_
timestamp 1676037725
transform 1 0 9108 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0587_
timestamp 1676037725
transform 1 0 26956 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0588_
timestamp 1676037725
transform 1 0 18216 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0589_
timestamp 1676037725
transform 1 0 27876 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1676037725
transform 1 0 23368 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0591_
timestamp 1676037725
transform 1 0 27324 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0592_
timestamp 1676037725
transform 1 0 21712 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0593_
timestamp 1676037725
transform 1 0 30360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0594_
timestamp 1676037725
transform 1 0 36064 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0595_
timestamp 1676037725
transform 1 0 24932 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0596_
timestamp 1676037725
transform 1 0 9108 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0597_
timestamp 1676037725
transform 1 0 9200 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0598_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0599_
timestamp 1676037725
transform 1 0 14996 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0600_
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0601_
timestamp 1676037725
transform 1 0 20148 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0602_
timestamp 1676037725
transform 1 0 14076 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0603_
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0604_
timestamp 1676037725
transform 1 0 16008 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1676037725
transform 1 0 25300 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0606_
timestamp 1676037725
transform 1 0 27968 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0607_
timestamp 1676037725
transform 1 0 28152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0608_
timestamp 1676037725
transform 1 0 19596 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0609_
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0610_
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_4  _0611_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34592 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0612_
timestamp 1676037725
transform 1 0 3956 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1676037725
transform 1 0 21068 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0614_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0615_
timestamp 1676037725
transform 1 0 32660 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0617_
timestamp 1676037725
transform 1 0 32292 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 1676037725
transform 1 0 30912 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 1676037725
transform 1 0 25116 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0620_
timestamp 1676037725
transform 1 0 28428 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0621_
timestamp 1676037725
transform 1 0 14996 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1676037725
transform 1 0 34408 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 1676037725
transform 1 0 24472 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0624_
timestamp 1676037725
transform 1 0 10028 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0625_
timestamp 1676037725
transform 1 0 32752 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1676037725
transform 1 0 30820 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0627_
timestamp 1676037725
transform 1 0 27508 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1676037725
transform 1 0 30728 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1676037725
transform 1 0 2300 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 1676037725
transform 1 0 2300 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0631_
timestamp 1676037725
transform 1 0 14904 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1676037725
transform 1 0 13616 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0633_
timestamp 1676037725
transform 1 0 20700 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1676037725
transform 1 0 23184 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 1676037725
transform 1 0 8832 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0637_
timestamp 1676037725
transform 1 0 26496 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0638_
timestamp 1676037725
transform 1 0 14444 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 1676037725
transform 1 0 32936 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0640_
timestamp 1676037725
transform 1 0 30360 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0641_
timestamp 1676037725
transform 1 0 12604 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1676037725
transform 1 0 12788 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0643_
timestamp 1676037725
transform 1 0 5428 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_2  _0644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34776 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0645_
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0646_
timestamp 1676037725
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0647_
timestamp 1676037725
transform 1 0 11408 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0648_
timestamp 1676037725
transform 1 0 26864 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0649_
timestamp 1676037725
transform 1 0 34960 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0650_
timestamp 1676037725
transform 1 0 24564 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0651_
timestamp 1676037725
transform 1 0 34868 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0652_
timestamp 1676037725
transform 1 0 10212 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0653_
timestamp 1676037725
transform 1 0 30176 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0654_
timestamp 1676037725
transform 1 0 17848 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0655_
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0656_
timestamp 1676037725
transform 1 0 17296 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0657_
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0658_
timestamp 1676037725
transform 1 0 37536 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0659_
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0660_
timestamp 1676037725
transform 1 0 12880 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0661_
timestamp 1676037725
transform 1 0 30452 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0662_
timestamp 1676037725
transform 1 0 7636 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0663_
timestamp 1676037725
transform 1 0 9384 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0664_
timestamp 1676037725
transform 1 0 12788 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0665_
timestamp 1676037725
transform 1 0 23000 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0666_
timestamp 1676037725
transform 1 0 11776 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0667_
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0668_
timestamp 1676037725
transform 1 0 5152 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0669_
timestamp 1676037725
transform 1 0 25760 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0670_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0671_
timestamp 1676037725
transform 1 0 34868 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1676037725
transform 1 0 27968 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0673_
timestamp 1676037725
transform 1 0 34868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0674_
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0675_
timestamp 1676037725
transform 1 0 36156 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0676_
timestamp 1676037725
transform 1 0 6624 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_4  _0677_
timestamp 1676037725
transform 1 0 35972 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0678_
timestamp 1676037725
transform 1 0 4324 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0679_
timestamp 1676037725
transform 1 0 19320 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0680_
timestamp 1676037725
transform 1 0 5244 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0681_
timestamp 1676037725
transform 1 0 33488 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0682_
timestamp 1676037725
transform 1 0 13340 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0683_
timestamp 1676037725
transform 1 0 33764 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 1676037725
transform 1 0 22356 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0685_
timestamp 1676037725
transform 1 0 4784 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0686_
timestamp 1676037725
transform 1 0 23184 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 1676037725
transform 1 0 2668 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0688_
timestamp 1676037725
transform 1 0 26128 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0689_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0691_
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0692_
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 1676037725
transform 1 0 25116 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0694_
timestamp 1676037725
transform 1 0 10396 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0697_
timestamp 1676037725
transform 1 0 14720 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1676037725
transform 1 0 30820 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1676037725
transform 1 0 18124 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0700_
timestamp 1676037725
transform 1 0 20056 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0701_
timestamp 1676037725
transform 1 0 4140 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 1676037725
transform 1 0 29440 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0703_
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1676037725
transform 1 0 20424 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1676037725
transform 1 0 29716 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0706_
timestamp 1676037725
transform 1 0 27784 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 1676037725
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0708_
timestamp 1676037725
transform 1 0 22172 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 1676037725
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_4  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__and2_1  _0711_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7544 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_4  _0712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_2  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10120 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_4  _0714_
timestamp 1676037725
transform 1 0 12420 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _0715_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2760 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _0717_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _0718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12420 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__and3_1  _0719_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0720_
timestamp 1676037725
transform 1 0 4416 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0721_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0722_
timestamp 1676037725
transform 1 0 34868 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0723_
timestamp 1676037725
transform 1 0 26036 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0724_
timestamp 1676037725
transform 1 0 34040 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0725_
timestamp 1676037725
transform 1 0 31648 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0726_
timestamp 1676037725
transform 1 0 28704 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0727_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0728_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0729_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0730_
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0731_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15824 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0732_
timestamp 1676037725
transform 1 0 30728 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0733_
timestamp 1676037725
transform 1 0 34868 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0734_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0735_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32752 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0736_
timestamp 1676037725
transform 1 0 27140 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0737_
timestamp 1676037725
transform 1 0 27140 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0738_
timestamp 1676037725
transform 1 0 29716 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0739_
timestamp 1676037725
transform 1 0 28152 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0740_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26956 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0741_
timestamp 1676037725
transform 1 0 26312 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1676037725
transform 1 0 25760 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0743_
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_2  _0744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26404 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0745_
timestamp 1676037725
transform 1 0 14628 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0746_
timestamp 1676037725
transform 1 0 17296 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0747_
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_2  _0748_
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0749_
timestamp 1676037725
transform 1 0 25576 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0750_
timestamp 1676037725
transform 1 0 27600 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0751_
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0752_
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0753_
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0754_
timestamp 1676037725
transform 1 0 6532 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0755_
timestamp 1676037725
transform 1 0 8004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0756_
timestamp 1676037725
transform 1 0 5612 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0757_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0758_
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0759_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0760_
timestamp 1676037725
transform 1 0 22908 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0761_
timestamp 1676037725
transform 1 0 21620 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0762_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0763_
timestamp 1676037725
transform 1 0 5428 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0764_
timestamp 1676037725
transform 1 0 6624 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0765_
timestamp 1676037725
transform 1 0 13248 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_4  _0766_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12328 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0767_
timestamp 1676037725
transform 1 0 19596 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0768_
timestamp 1676037725
transform 1 0 14720 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0769_
timestamp 1676037725
transform 1 0 19872 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0770_
timestamp 1676037725
transform 1 0 20608 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0771_
timestamp 1676037725
transform 1 0 13156 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0772_
timestamp 1676037725
transform 1 0 14904 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0773_
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_2  _0774_
timestamp 1676037725
transform 1 0 14628 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0775_
timestamp 1676037725
transform 1 0 10120 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0776_
timestamp 1676037725
transform 1 0 9016 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0777_
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_4  _0778_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _0779_
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0780_
timestamp 1676037725
transform 1 0 2760 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0781_
timestamp 1676037725
transform 1 0 1840 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0782_
timestamp 1676037725
transform 1 0 4048 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0783_
timestamp 1676037725
transform 1 0 5244 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0784_
timestamp 1676037725
transform 1 0 22724 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0785_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0786_
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0787_
timestamp 1676037725
transform 1 0 22356 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0788_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0789_
timestamp 1676037725
transform 1 0 2024 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0790_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0791_
timestamp 1676037725
transform 1 0 3956 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0792_
timestamp 1676037725
transform 1 0 13156 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0793_
timestamp 1676037725
transform 1 0 1656 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0794_
timestamp 1676037725
transform 1 0 28704 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0795_
timestamp 1676037725
transform 1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0796_
timestamp 1676037725
transform 1 0 32384 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0797_
timestamp 1676037725
transform 1 0 31372 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0798_
timestamp 1676037725
transform 1 0 31556 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0799_
timestamp 1676037725
transform 1 0 27324 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0800_
timestamp 1676037725
transform 1 0 25944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0801_
timestamp 1676037725
transform 1 0 33672 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0802_
timestamp 1676037725
transform 1 0 33580 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0803_
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0804_
timestamp 1676037725
transform 1 0 17204 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0805_
timestamp 1676037725
transform 1 0 12880 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0806_
timestamp 1676037725
transform 1 0 8096 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_2  _0807_
timestamp 1676037725
transform 1 0 15916 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0808_
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0809_
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0810_
timestamp 1676037725
transform 1 0 10396 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0811_
timestamp 1676037725
transform 1 0 18308 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0812_
timestamp 1676037725
transform 1 0 18124 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0813_
timestamp 1676037725
transform 1 0 28704 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0814_
timestamp 1676037725
transform 1 0 32752 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0815_
timestamp 1676037725
transform 1 0 29440 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_2  _0816_
timestamp 1676037725
transform 1 0 30360 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0817_
timestamp 1676037725
transform 1 0 17480 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0818_
timestamp 1676037725
transform 1 0 17112 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0819_
timestamp 1676037725
transform 1 0 6808 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0820_
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0821_
timestamp 1676037725
transform 1 0 11684 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0822_
timestamp 1676037725
transform 1 0 26588 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0823_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0824_
timestamp 1676037725
transform 1 0 31648 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0825_
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0826_
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0827_
timestamp 1676037725
transform 1 0 5612 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0828_
timestamp 1676037725
transform 1 0 5428 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0829_
timestamp 1676037725
transform 1 0 4508 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0830_
timestamp 1676037725
transform 1 0 14352 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0831_
timestamp 1676037725
transform 1 0 5704 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0832_
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0833_
timestamp 1676037725
transform 1 0 32384 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0834_
timestamp 1676037725
transform 1 0 30820 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0835_
timestamp 1676037725
transform 1 0 32476 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0836_
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0837_
timestamp 1676037725
transform 1 0 33488 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0838_
timestamp 1676037725
transform 1 0 25760 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_2  _0839_
timestamp 1676037725
transform 1 0 25760 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0840_
timestamp 1676037725
transform 1 0 16928 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0841_
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0842_
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0843_
timestamp 1676037725
transform 1 0 25760 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0844_
timestamp 1676037725
transform 1 0 35972 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0845_
timestamp 1676037725
transform 1 0 33580 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0846_
timestamp 1676037725
transform 1 0 24656 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0847_
timestamp 1676037725
transform 1 0 33396 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0848_
timestamp 1676037725
transform 1 0 35052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0849_
timestamp 1676037725
transform 1 0 11960 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0850_
timestamp 1676037725
transform 1 0 3956 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0851_
timestamp 1676037725
transform 1 0 12328 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0852_
timestamp 1676037725
transform 1 0 10396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0853_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0854_
timestamp 1676037725
transform 1 0 20884 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0855_
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0857_
timestamp 1676037725
transform 1 0 22080 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0858_
timestamp 1676037725
transform 1 0 10948 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0859_
timestamp 1676037725
transform 1 0 7728 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0860_
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0861_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0862_
timestamp 1676037725
transform 1 0 7544 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1676037725
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1676037725
transform 1 0 13984 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1676037725
transform 1 0 37168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1676037725
transform 1 0 4508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1676037725
transform 1 0 36064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1676037725
transform 1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1676037725
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1676037725
transform 1 0 37444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1676037725
transform 1 0 33764 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1676037725
transform 1 0 13156 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1676037725
transform 1 0 37168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1676037725
transform 1 0 33856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1676037725
transform 1 0 36524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1676037725
transform 1 0 30544 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1676037725
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1676037725
transform 1 0 13984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1676037725
transform 1 0 35880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1676037725
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1676037725
transform 1 0 36708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1676037725
transform 1 0 6164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1676037725
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1676037725
transform 1 0 8096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1676037725
transform 1 0 38456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1676037725
transform 1 0 26312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1676037725
transform 1 0 36800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1676037725
transform 1 0 36708 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1676037725
transform 1 0 37904 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1676037725
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1676037725
transform 1 0 6808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1676037725
transform 1 0 9016 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1676037725
transform 1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1676037725
transform 1 0 38364 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1676037725
transform 1 0 34040 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1676037725
transform 1 0 36616 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0913_
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1676037725
transform 1 0 18584 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0915_
timestamp 1676037725
transform 1 0 37168 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1676037725
transform 1 0 28060 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1676037725
transform 1 0 31004 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1676037725
transform 1 0 5612 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1676037725
transform 1 0 37536 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1676037725
transform 1 0 29716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1676037725
transform 1 0 38088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1676037725
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1676037725
transform 1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1676037725
transform 1 0 10304 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1676037725
transform 1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1676037725
transform 1 0 16100 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1676037725
transform 1 0 37536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1676037725
transform 1 0 38180 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1676037725
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0932_
timestamp 1676037725
transform 1 0 30084 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1676037725
transform 1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1676037725
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1676037725
transform 1 0 37536 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1676037725
transform 1 0 38088 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1676037725
transform 1 0 2576 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1676037725
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1676037725
transform 1 0 28520 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1676037725
transform 1 0 28152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1676037725
transform 1 0 38088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0945_
timestamp 1676037725
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1676037725
transform 1 0 31556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1676037725
transform 1 0 36156 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1676037725
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1676037725
transform 1 0 27784 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1676037725
transform 1 0 31556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1676037725
transform 1 0 28612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1676037725
transform 1 0 35512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1676037725
transform 1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1676037725
transform 1 0 37996 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1676037725
transform 1 0 23920 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1676037725
transform 1 0 5520 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1676037725
transform 1 0 34132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1676037725
transform 1 0 9660 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1676037725
transform 1 0 12972 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1676037725
transform 1 0 36708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1676037725
transform 1 0 38088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1676037725
transform 1 0 36064 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1676037725
transform 1 0 15824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1676037725
transform 1 0 37720 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1676037725
transform 1 0 17848 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1676037725
transform 1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1676037725
transform 1 0 36708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1676037725
transform 1 0 38456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1676037725
transform 1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1676037725
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1676037725
transform 1 0 29716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1676037725
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0981_
timestamp 1676037725
transform 1 0 16836 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1676037725
transform 1 0 5152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1676037725
transform 1 0 23828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1676037725
transform 1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1676037725
transform 1 0 34132 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1676037725
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1676037725
transform 1 0 2576 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1676037725
transform 1 0 35696 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0992_
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0993_
timestamp 1676037725
transform 1 0 29164 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1676037725
transform 1 0 4324 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1676037725
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1676037725
transform 1 0 34132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1676037725
transform 1 0 11776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1676037725
transform 1 0 28520 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1676037725
transform 1 0 10304 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1676037725
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1676037725
transform 1 0 2668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1676037725
transform 1 0 2668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1676037725
transform 1 0 34592 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1676037725
transform 1 0 26404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1676037725
transform 1 0 2576 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1676037725
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1676037725
transform 1 0 31280 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1676037725
transform 1 0 6256 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1676037725
transform 1 0 37352 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1676037725
transform 1 0 4968 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1676037725
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1676037725
transform 1 0 21252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1676037725
transform 1 0 33764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1021_
timestamp 1676037725
transform 1 0 2024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1676037725
transform 1 0 38088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1676037725
transform 1 0 2852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1676037725
transform 1 0 16468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1676037725
transform 1 0 37812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1676037725
transform 1 0 37444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1676037725
transform 1 0 6164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1676037725
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1676037725
transform 1 0 30176 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1676037725
transform 1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1676037725
transform 1 0 36064 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1676037725
transform 1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1676037725
transform 1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1676037725
transform 1 0 6256 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1676037725
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1676037725
transform 1 0 2208 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1676037725
transform 1 0 37536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1676037725
transform 1 0 37812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1676037725
transform 1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1676037725
transform 1 0 9660 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1676037725
transform 1 0 31832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1676037725
transform 1 0 12052 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1676037725
transform 1 0 6164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1676037725
transform 1 0 23644 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1676037725
transform 1 0 37444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1676037725
transform 1 0 31924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1676037725
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1676037725
transform 1 0 32476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1676037725
transform 1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1055_
timestamp 1676037725
transform 1 0 24840 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1056_
timestamp 1676037725
transform 1 0 13248 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1057_
timestamp 1676037725
transform 1 0 26864 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1058_
timestamp 1676037725
transform 1 0 28152 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1060_
timestamp 1676037725
transform 1 0 2208 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26772 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1062_
timestamp 1676037725
transform 1 0 2392 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1063_
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1064_
timestamp 1676037725
transform 1 0 14904 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1065_
timestamp 1676037725
transform 1 0 31004 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1066_
timestamp 1676037725
transform 1 0 13156 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1067_
timestamp 1676037725
transform 1 0 12420 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1068_
timestamp 1676037725
transform 1 0 6164 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1069_
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1070_
timestamp 1676037725
transform 1 0 27232 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1071_
timestamp 1676037725
transform 1 0 15272 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1072_
timestamp 1676037725
transform 1 0 34960 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1073_
timestamp 1676037725
transform 1 0 2668 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1074_
timestamp 1676037725
transform 1 0 13892 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1075_
timestamp 1676037725
transform 1 0 24840 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1076_
timestamp 1676037725
transform 1 0 1656 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1077_
timestamp 1676037725
transform 1 0 20608 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1078_
timestamp 1676037725
transform 1 0 2760 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1079_
timestamp 1676037725
transform 1 0 22264 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1080_
timestamp 1676037725
transform 1 0 27416 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1081_
timestamp 1676037725
transform 1 0 19044 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1082_
timestamp 1676037725
transform 1 0 33120 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1083_
timestamp 1676037725
transform 1 0 6808 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1084_
timestamp 1676037725
transform 1 0 18216 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1085_
timestamp 1676037725
transform 1 0 2576 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1086_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1087_
timestamp 1676037725
transform 1 0 32568 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1088_
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1089_
timestamp 1676037725
transform 1 0 34868 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1090_
timestamp 1676037725
transform 1 0 24748 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1091_
timestamp 1676037725
transform 1 0 24196 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1092_
timestamp 1676037725
transform 1 0 24564 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1093_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1094_
timestamp 1676037725
transform 1 0 25024 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1095_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1096_
timestamp 1676037725
transform 1 0 11316 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1097_
timestamp 1676037725
transform 1 0 20976 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1098_
timestamp 1676037725
transform 1 0 11040 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1099_
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1100_
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1101_
timestamp 1676037725
transform 1 0 30728 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1676037725
transform 1 0 10672 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 1676037725
transform 1 0 35144 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1104_
timestamp 1676037725
transform 1 0 35052 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1105_
timestamp 1676037725
transform 1 0 5152 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 1676037725
transform 1 0 17112 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1107_
timestamp 1676037725
transform 1 0 1748 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 1676037725
transform 1 0 15364 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 1676037725
transform 1 0 29624 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1111_
timestamp 1676037725
transform 1 0 32292 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1113_
timestamp 1676037725
transform 1 0 35880 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1114_
timestamp 1676037725
transform 1 0 9568 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1115_
timestamp 1676037725
transform 1 0 11684 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1116_
timestamp 1676037725
transform 1 0 20792 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1117_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1118_
timestamp 1676037725
transform 1 0 34868 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1119_
timestamp 1676037725
transform 1 0 14260 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1676037725
transform 1 0 16928 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1121_
timestamp 1676037725
transform 1 0 22632 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 1676037725
transform 1 0 30544 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 1676037725
transform 1 0 14536 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1124_
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1126_
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1127_
timestamp 1676037725
transform 1 0 32292 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 1676037725
transform 1 0 11960 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1131_
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1132_
timestamp 1676037725
transform 1 0 2852 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1133_
timestamp 1676037725
transform 1 0 31004 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1134_
timestamp 1676037725
transform 1 0 27140 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1676037725
transform 1 0 25116 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 1676037725
transform 1 0 34868 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1137_
timestamp 1676037725
transform 1 0 35052 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 1676037725
transform 1 0 22264 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1139_
timestamp 1676037725
transform 1 0 30176 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1140_
timestamp 1676037725
transform 1 0 20608 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1141_
timestamp 1676037725
transform 1 0 28152 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1142_
timestamp 1676037725
transform 1 0 25116 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1143_
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1144_
timestamp 1676037725
transform 1 0 32292 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1145_
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1146_
timestamp 1676037725
transform 1 0 34868 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1147_
timestamp 1676037725
transform 1 0 10764 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1148_
timestamp 1676037725
transform 1 0 20792 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1149_
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1150_
timestamp 1676037725
transform 1 0 6256 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1151_
timestamp 1676037725
transform 1 0 29716 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1152_
timestamp 1676037725
transform 1 0 28612 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1153_
timestamp 1676037725
transform 1 0 12696 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1154_
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1155_
timestamp 1676037725
transform 1 0 12880 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1156_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1157_
timestamp 1676037725
transform 1 0 29716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1676037725
transform 1 0 10580 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 1676037725
transform 1 0 22172 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1160_
timestamp 1676037725
transform 1 0 28612 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1161_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 1676037725
transform 1 0 15916 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1163_
timestamp 1676037725
transform 1 0 6532 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1164_
timestamp 1676037725
transform 1 0 7084 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1165_
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1166_
timestamp 1676037725
transform 1 0 32292 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1676037725
transform 1 0 29440 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1676037725
transform 1 0 23092 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1169_
timestamp 1676037725
transform 1 0 19044 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1170_
timestamp 1676037725
transform 1 0 23092 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1676037725
transform 1 0 14352 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1173_
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1174_
timestamp 1676037725
transform 1 0 8280 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1175_
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1676037725
transform 1 0 22356 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1676037725
transform 1 0 19320 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1178_
timestamp 1676037725
transform 1 0 34592 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1179_
timestamp 1676037725
transform 1 0 27324 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 1676037725
transform 1 0 19320 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1183_
timestamp 1676037725
transform 1 0 24748 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1184_
timestamp 1676037725
transform 1 0 34868 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1185_
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1187_
timestamp 1676037725
transform 1 0 2392 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1188_
timestamp 1676037725
transform 1 0 15916 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1189_
timestamp 1676037725
transform 1 0 11960 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1190_
timestamp 1676037725
transform 1 0 35972 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1676037725
transform 1 0 28244 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1192_
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1193_
timestamp 1676037725
transform 1 0 10764 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1194_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1195_
timestamp 1676037725
transform 1 0 15456 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 1676037725
transform 1 0 14536 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1197_
timestamp 1676037725
transform 1 0 20516 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1676037725
transform 1 0 2944 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1199_
timestamp 1676037725
transform 1 0 33120 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1200_
timestamp 1676037725
transform 1 0 27140 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1201_
timestamp 1676037725
transform 1 0 2300 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1202_
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1203_
timestamp 1676037725
transform 1 0 30544 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1204_
timestamp 1676037725
transform 1 0 7544 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1205_
timestamp 1676037725
transform 1 0 36800 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1206_
timestamp 1676037725
transform 1 0 5888 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1676037725
transform 1 0 34500 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1208_
timestamp 1676037725
transform 1 0 13892 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1210_
timestamp 1676037725
transform 1 0 32568 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 1676037725
transform 1 0 3680 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1676037725
transform 1 0 25668 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1213_
timestamp 1676037725
transform 1 0 36800 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1214_
timestamp 1676037725
transform 1 0 4232 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1215_
timestamp 1676037725
transform 1 0 31924 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1216_
timestamp 1676037725
transform 1 0 2208 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1217_
timestamp 1676037725
transform 1 0 19504 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1218_
timestamp 1676037725
transform 1 0 32016 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1676037725
transform 1 0 29992 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 1676037725
transform 1 0 9752 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1221_
timestamp 1676037725
transform 1 0 23736 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1222_
timestamp 1676037725
transform 1 0 16744 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1223_
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1224_
timestamp 1676037725
transform 1 0 17940 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1225_
timestamp 1676037725
transform 1 0 34868 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1226_
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1227_
timestamp 1676037725
transform 1 0 19320 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1228_
timestamp 1676037725
transform 1 0 4600 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1229_
timestamp 1676037725
transform 1 0 19780 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1230_
timestamp 1676037725
transform 1 0 3956 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1231_
timestamp 1676037725
transform 1 0 29716 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1232_
timestamp 1676037725
transform 1 0 20424 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1233_
timestamp 1676037725
transform 1 0 5888 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1234_
timestamp 1676037725
transform 1 0 2208 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1235_
timestamp 1676037725
transform 1 0 28796 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1236_
timestamp 1676037725
transform 1 0 4968 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1237_
timestamp 1676037725
transform 1 0 31280 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1238_
timestamp 1676037725
transform 1 0 7636 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1239_
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1240_
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1241_
timestamp 1676037725
transform 1 0 29624 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1242_
timestamp 1676037725
transform 1 0 15640 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1243_
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1244_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1245_
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7636 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1676037725
transform 1 0 9292 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1676037725
transform 1 0 14904 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1676037725
transform 1 0 14904 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1676037725
transform 1 0 7176 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1676037725
transform 1 0 6900 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1676037725
transform 1 0 25484 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1676037725
transform 1 0 32660 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1676037725
transform 1 0 32660 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1676037725
transform 1 0 31372 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1676037725
transform 1 0 30820 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout73 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18400 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout74 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12328 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout75
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout77
timestamp 1676037725
transform 1 0 8740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout78
timestamp 1676037725
transform 1 0 12880 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout79
timestamp 1676037725
transform 1 0 22448 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 1676037725
transform 1 0 21160 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout82
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout83
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout84
timestamp 1676037725
transform 1 0 14720 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout85
timestamp 1676037725
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout86
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout87
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout88
timestamp 1676037725
transform 1 0 9476 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout89
timestamp 1676037725
transform 1 0 9200 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout90
timestamp 1676037725
transform 1 0 18400 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout91
timestamp 1676037725
transform 1 0 22632 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout92
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout93
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout94
timestamp 1676037725
transform 1 0 20240 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout95
timestamp 1676037725
transform 1 0 20148 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout96
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout97
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout98
timestamp 1676037725
transform 1 0 17204 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout99
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout100 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14628 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout101
timestamp 1676037725
transform 1 0 12972 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout102
timestamp 1676037725
transform 1 0 35328 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout103
timestamp 1676037725
transform 1 0 34960 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout104
timestamp 1676037725
transform 1 0 12420 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout105
timestamp 1676037725
transform 1 0 34776 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout106
timestamp 1676037725
transform 1 0 35604 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout107
timestamp 1676037725
transform 1 0 35604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout108
timestamp 1676037725
transform 1 0 11684 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout109
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout110
timestamp 1676037725
transform 1 0 35604 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout111
timestamp 1676037725
transform 1 0 31188 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout112
timestamp 1676037725
transform 1 0 18492 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout113
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout114
timestamp 1676037725
transform 1 0 27416 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout115
timestamp 1676037725
transform 1 0 37076 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout116
timestamp 1676037725
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout117
timestamp 1676037725
transform 1 0 17848 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout118
timestamp 1676037725
transform 1 0 33304 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout119
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout120
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout121
timestamp 1676037725
transform 1 0 9016 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout122
timestamp 1676037725
transform 1 0 32476 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout123
timestamp 1676037725
transform 1 0 32568 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout124
timestamp 1676037725
transform 1 0 7820 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout125
timestamp 1676037725
transform 1 0 9476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout126
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout127
timestamp 1676037725
transform 1 0 17020 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout128
timestamp 1676037725
transform 1 0 12972 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout129
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout130
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout131
timestamp 1676037725
transform 1 0 4968 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout132
timestamp 1676037725
transform 1 0 3864 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout133
timestamp 1676037725
transform 1 0 15272 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout134
timestamp 1676037725
transform 1 0 18308 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout135
timestamp 1676037725
transform 1 0 23092 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout136
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout137
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout138
timestamp 1676037725
transform 1 0 24564 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout139
timestamp 1676037725
transform 1 0 23184 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout140
timestamp 1676037725
transform 1 0 30912 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout141
timestamp 1676037725
transform 1 0 33948 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout142
timestamp 1676037725
transform 1 0 35512 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout143
timestamp 1676037725
transform 1 0 34868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout144
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout145
timestamp 1676037725
transform 1 0 23552 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout146
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout147
timestamp 1676037725
transform 1 0 29716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout148
timestamp 1676037725
transform 1 0 29348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout149
timestamp 1676037725
transform 1 0 22540 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout150
timestamp 1676037725
transform 1 0 11500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  fanout151 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout152
timestamp 1676037725
transform 1 0 10580 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  fanout153
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout154
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1676037725
transform 1 0 29716 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1676037725
transform 1 0 11684 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1676037725
transform 1 0 23184 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1676037725
transform 1 0 6532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1676037725
transform 1 0 21988 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1676037725
transform 1 0 18124 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 1676037725
transform 1 0 25208 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input12
timestamp 1676037725
transform 1 0 3956 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input14
timestamp 1676037725
transform 1 0 1564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input15
timestamp 1676037725
transform 1 0 23276 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 1676037725
transform 1 0 30636 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1676037725
transform 1 0 38180 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input19
timestamp 1676037725
transform 1 0 1564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1676037725
transform 1 0 38180 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input22
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input23
timestamp 1676037725
transform 1 0 13248 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input24
timestamp 1676037725
transform 1 0 37904 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input25
timestamp 1676037725
transform 1 0 35328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1676037725
transform 1 0 12972 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input27
timestamp 1676037725
transform 1 0 38180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input28
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input29
timestamp 1676037725
transform 1 0 2024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 1676037725
transform 1 0 38180 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input32
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1676037725
transform 1 0 36156 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1676037725
transform 1 0 34868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input35
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input36
timestamp 1676037725
transform 1 0 14904 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input37
timestamp 1676037725
transform 1 0 20976 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input39
timestamp 1676037725
transform 1 0 2024 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 1676037725
transform 1 0 38364 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output41
timestamp 1676037725
transform 1 0 3128 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output42
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output43
timestamp 1676037725
transform 1 0 27140 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output44
timestamp 1676037725
transform 1 0 7820 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output45
timestamp 1676037725
transform 1 0 37444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output46
timestamp 1676037725
transform 1 0 2944 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output47
timestamp 1676037725
transform 1 0 33304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output48
timestamp 1676037725
transform 1 0 1564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output49
timestamp 1676037725
transform 1 0 38364 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output50
timestamp 1676037725
transform 1 0 38364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output51
timestamp 1676037725
transform 1 0 20056 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output52
timestamp 1676037725
transform 1 0 29716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output53
timestamp 1676037725
transform 1 0 38364 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output54
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output55
timestamp 1676037725
transform 1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output56
timestamp 1676037725
transform 1 0 32292 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output57
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output58
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output59
timestamp 1676037725
transform 1 0 38364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1676037725
transform 1 0 32292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1676037725
transform 1 0 16836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1676037725
transform 1 0 10856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1676037725
transform 1 0 28888 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1676037725
transform 1 0 36432 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 28998 28354 29054 29154 0 FreeSans 224 90 0 0 read_address[0]
port 1 nsew signal input
flabel metal2 s 10966 28354 11022 29154 0 FreeSans 224 90 0 0 read_address[1]
port 2 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 read_address[2]
port 3 nsew signal input
flabel metal3 s 39566 18368 40366 18488 0 FreeSans 480 0 0 0 read_address[3]
port 4 nsew signal input
flabel metal3 s 39566 22448 40366 22568 0 FreeSans 480 0 0 0 read_address[4]
port 5 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 read_data[0]
port 6 nsew signal tristate
flabel metal3 s 39566 2048 40366 2168 0 FreeSans 480 0 0 0 read_data[10]
port 7 nsew signal tristate
flabel metal2 s 27066 28354 27122 29154 0 FreeSans 224 90 0 0 read_data[11]
port 8 nsew signal tristate
flabel metal2 s 7746 28354 7802 29154 0 FreeSans 224 90 0 0 read_data[12]
port 9 nsew signal tristate
flabel metal2 s 37370 28354 37426 29154 0 FreeSans 224 90 0 0 read_data[13]
port 10 nsew signal tristate
flabel metal2 s 662 28354 718 29154 0 FreeSans 224 90 0 0 read_data[14]
port 11 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 read_data[15]
port 12 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 read_data[16]
port 13 nsew signal tristate
flabel metal3 s 39566 7488 40366 7608 0 FreeSans 480 0 0 0 read_data[17]
port 14 nsew signal tristate
flabel metal3 s 39566 3408 40366 3528 0 FreeSans 480 0 0 0 read_data[18]
port 15 nsew signal tristate
flabel metal2 s 19982 28354 20038 29154 0 FreeSans 224 90 0 0 read_data[19]
port 16 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 read_data[1]
port 17 nsew signal tristate
flabel metal2 s 39302 28354 39358 29154 0 FreeSans 224 90 0 0 read_data[20]
port 18 nsew signal tristate
flabel metal3 s 39566 8 40366 128 0 FreeSans 480 0 0 0 read_data[21]
port 19 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 read_data[22]
port 20 nsew signal tristate
flabel metal2 s 32218 28354 32274 29154 0 FreeSans 224 90 0 0 read_data[23]
port 21 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 read_data[24]
port 22 nsew signal tristate
flabel metal3 s 39566 17008 40366 17128 0 FreeSans 480 0 0 0 read_data[25]
port 23 nsew signal tristate
flabel metal3 s 39566 20408 40366 20528 0 FreeSans 480 0 0 0 read_data[26]
port 24 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 read_data[27]
port 25 nsew signal tristate
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 read_data[28]
port 26 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 read_data[29]
port 27 nsew signal tristate
flabel metal2 s 16118 28354 16174 29154 0 FreeSans 224 90 0 0 read_data[2]
port 28 nsew signal tristate
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 read_data[30]
port 29 nsew signal tristate
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 read_data[31]
port 30 nsew signal tristate
flabel metal3 s 39566 14968 40366 15088 0 FreeSans 480 0 0 0 read_data[3]
port 31 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 read_data[4]
port 32 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 read_data[5]
port 33 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 read_data[6]
port 34 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 read_data[7]
port 35 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 read_data[8]
port 36 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 read_data[9]
port 37 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 reset
port 38 nsew signal input
flabel metal4 s 5705 2128 6025 26704 0 FreeSans 1920 90 0 0 vccd1
port 39 nsew power bidirectional
flabel metal4 s 15227 2128 15547 26704 0 FreeSans 1920 90 0 0 vccd1
port 39 nsew power bidirectional
flabel metal4 s 24749 2128 25069 26704 0 FreeSans 1920 90 0 0 vccd1
port 39 nsew power bidirectional
flabel metal4 s 34271 2128 34591 26704 0 FreeSans 1920 90 0 0 vccd1
port 39 nsew power bidirectional
flabel metal4 s 10466 2128 10786 26704 0 FreeSans 1920 90 0 0 vssd1
port 40 nsew ground bidirectional
flabel metal4 s 19988 2128 20308 26704 0 FreeSans 1920 90 0 0 vssd1
port 40 nsew ground bidirectional
flabel metal4 s 29510 2128 29830 26704 0 FreeSans 1920 90 0 0 vssd1
port 40 nsew ground bidirectional
flabel metal4 s 39032 2128 39352 26704 0 FreeSans 1920 90 0 0 vssd1
port 40 nsew ground bidirectional
flabel metal2 s 5814 28354 5870 29154 0 FreeSans 224 90 0 0 write_address[0]
port 41 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 write_address[1]
port 42 nsew signal input
flabel metal2 s 21914 28354 21970 29154 0 FreeSans 224 90 0 0 write_address[2]
port 43 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 write_address[3]
port 44 nsew signal input
flabel metal3 s 39566 5448 40366 5568 0 FreeSans 480 0 0 0 write_address[4]
port 45 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 write_data[0]
port 46 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 write_data[10]
port 47 nsew signal input
flabel metal2 s 18050 28354 18106 29154 0 FreeSans 224 90 0 0 write_data[11]
port 48 nsew signal input
flabel metal2 s 25134 28354 25190 29154 0 FreeSans 224 90 0 0 write_data[12]
port 49 nsew signal input
flabel metal2 s 3882 28354 3938 29154 0 FreeSans 224 90 0 0 write_data[13]
port 50 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 write_data[14]
port 51 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 write_data[15]
port 52 nsew signal input
flabel metal2 s 23202 28354 23258 29154 0 FreeSans 224 90 0 0 write_data[16]
port 53 nsew signal input
flabel metal2 s 30286 28354 30342 29154 0 FreeSans 224 90 0 0 write_data[17]
port 54 nsew signal input
flabel metal3 s 39566 27888 40366 28008 0 FreeSans 480 0 0 0 write_data[18]
port 55 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 write_data[19]
port 56 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 write_data[1]
port 57 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 write_data[20]
port 58 nsew signal input
flabel metal3 s 39566 25848 40366 25968 0 FreeSans 480 0 0 0 write_data[21]
port 59 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 write_data[22]
port 60 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 write_data[23]
port 61 nsew signal input
flabel metal3 s 39566 24488 40366 24608 0 FreeSans 480 0 0 0 write_data[24]
port 62 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 write_data[25]
port 63 nsew signal input
flabel metal2 s 12898 28354 12954 29154 0 FreeSans 224 90 0 0 write_data[26]
port 64 nsew signal input
flabel metal3 s 39566 10888 40366 11008 0 FreeSans 480 0 0 0 write_data[27]
port 65 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 write_data[28]
port 66 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 write_data[29]
port 67 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 write_data[2]
port 68 nsew signal input
flabel metal3 s 39566 12928 40366 13048 0 FreeSans 480 0 0 0 write_data[30]
port 69 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 write_data[31]
port 70 nsew signal input
flabel metal2 s 36082 28354 36138 29154 0 FreeSans 224 90 0 0 write_data[3]
port 71 nsew signal input
flabel metal2 s 34150 28354 34206 29154 0 FreeSans 224 90 0 0 write_data[4]
port 72 nsew signal input
flabel metal2 s 9034 28354 9090 29154 0 FreeSans 224 90 0 0 write_data[5]
port 73 nsew signal input
flabel metal2 s 14830 28354 14886 29154 0 FreeSans 224 90 0 0 write_data[6]
port 74 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 write_data[7]
port 75 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 write_data[8]
port 76 nsew signal input
flabel metal2 s 1950 28354 2006 29154 0 FreeSans 224 90 0 0 write_data[9]
port 77 nsew signal input
flabel metal3 s 39566 9528 40366 9648 0 FreeSans 480 0 0 0 write_enable
port 78 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40366 29154
<< end >>
