VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Scalar_Register_File
  CLASS BLOCK ;
  FOREIGN Scalar_Register_File ;
  ORIGIN 0.000 0.000 ;
  SIZE 201.830 BY 145.770 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END clk
  PIN read_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 141.770 145.270 145.770 ;
    END
  END read_address[0]
  PIN read_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 141.770 55.110 145.770 ;
    END
  END read_address[1]
  PIN read_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END read_address[2]
  PIN read_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 91.840 201.830 92.440 ;
    END
  END read_address[3]
  PIN read_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 112.240 201.830 112.840 ;
    END
  END read_address[4]
  PIN read_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END read_data[0]
  PIN read_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 10.240 201.830 10.840 ;
    END
  END read_data[10]
  PIN read_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 141.770 135.610 145.770 ;
    END
  END read_data[11]
  PIN read_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 141.770 39.010 145.770 ;
    END
  END read_data[12]
  PIN read_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 141.770 187.130 145.770 ;
    END
  END read_data[13]
  PIN read_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 141.770 3.590 145.770 ;
    END
  END read_data[14]
  PIN read_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END read_data[15]
  PIN read_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END read_data[16]
  PIN read_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 37.440 201.830 38.040 ;
    END
  END read_data[17]
  PIN read_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 17.040 201.830 17.640 ;
    END
  END read_data[18]
  PIN read_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 141.770 100.190 145.770 ;
    END
  END read_data[19]
  PIN read_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END read_data[1]
  PIN read_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 141.770 196.790 145.770 ;
    END
  END read_data[20]
  PIN read_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 0.040 201.830 0.640 ;
    END
  END read_data[21]
  PIN read_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END read_data[22]
  PIN read_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 141.770 161.370 145.770 ;
    END
  END read_data[23]
  PIN read_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END read_data[24]
  PIN read_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 85.040 201.830 85.640 ;
    END
  END read_data[25]
  PIN read_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 102.040 201.830 102.640 ;
    END
  END read_data[26]
  PIN read_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END read_data[27]
  PIN read_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END read_data[28]
  PIN read_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END read_data[29]
  PIN read_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 141.770 80.870 145.770 ;
    END
  END read_data[2]
  PIN read_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END read_data[30]
  PIN read_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END read_data[31]
  PIN read_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 74.840 201.830 75.440 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END read_data[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.525 10.640 30.125 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.135 10.640 77.735 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.745 10.640 125.345 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.355 10.640 172.955 133.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 52.330 10.640 53.930 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.940 10.640 101.540 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 147.550 10.640 149.150 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 195.160 10.640 196.760 133.520 ;
    END
  END vssd1
  PIN write_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 141.770 29.350 145.770 ;
    END
  END write_address[0]
  PIN write_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END write_address[1]
  PIN write_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 141.770 109.850 145.770 ;
    END
  END write_address[2]
  PIN write_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END write_address[3]
  PIN write_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 27.240 201.830 27.840 ;
    END
  END write_address[4]
  PIN write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END write_data[0]
  PIN write_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END write_data[10]
  PIN write_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 141.770 90.530 145.770 ;
    END
  END write_data[11]
  PIN write_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 141.770 125.950 145.770 ;
    END
  END write_data[12]
  PIN write_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 141.770 19.690 145.770 ;
    END
  END write_data[13]
  PIN write_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END write_data[14]
  PIN write_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END write_data[15]
  PIN write_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 141.770 116.290 145.770 ;
    END
  END write_data[16]
  PIN write_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 141.770 151.710 145.770 ;
    END
  END write_data[17]
  PIN write_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 139.440 201.830 140.040 ;
    END
  END write_data[18]
  PIN write_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END write_data[19]
  PIN write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END write_data[1]
  PIN write_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END write_data[20]
  PIN write_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 129.240 201.830 129.840 ;
    END
  END write_data[21]
  PIN write_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END write_data[22]
  PIN write_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END write_data[23]
  PIN write_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 122.440 201.830 123.040 ;
    END
  END write_data[24]
  PIN write_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END write_data[25]
  PIN write_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 141.770 64.770 145.770 ;
    END
  END write_data[26]
  PIN write_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 54.440 201.830 55.040 ;
    END
  END write_data[27]
  PIN write_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END write_data[28]
  PIN write_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END write_data[29]
  PIN write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END write_data[2]
  PIN write_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 64.640 201.830 65.240 ;
    END
  END write_data[30]
  PIN write_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END write_data[31]
  PIN write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 141.770 180.690 145.770 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 141.770 171.030 145.770 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 141.770 45.450 145.770 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 141.770 74.430 145.770 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 141.770 10.030 145.770 ;
    END
  END write_data[9]
  PIN write_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.830 47.640 201.830 48.240 ;
    END
  END write_enable
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 195.960 133.365 ;
      LAYER met1 ;
        RECT 0.070 0.380 197.730 141.400 ;
      LAYER met2 ;
        RECT 0.100 141.490 3.030 142.530 ;
        RECT 3.870 141.490 9.470 142.530 ;
        RECT 10.310 141.490 19.130 142.530 ;
        RECT 19.970 141.490 28.790 142.530 ;
        RECT 29.630 141.490 38.450 142.530 ;
        RECT 39.290 141.490 44.890 142.530 ;
        RECT 45.730 141.490 54.550 142.530 ;
        RECT 55.390 141.490 64.210 142.530 ;
        RECT 65.050 141.490 73.870 142.530 ;
        RECT 74.710 141.490 80.310 142.530 ;
        RECT 81.150 141.490 89.970 142.530 ;
        RECT 90.810 141.490 99.630 142.530 ;
        RECT 100.470 141.490 109.290 142.530 ;
        RECT 110.130 141.490 115.730 142.530 ;
        RECT 116.570 141.490 125.390 142.530 ;
        RECT 126.230 141.490 135.050 142.530 ;
        RECT 135.890 141.490 144.710 142.530 ;
        RECT 145.550 141.490 151.150 142.530 ;
        RECT 151.990 141.490 160.810 142.530 ;
        RECT 161.650 141.490 170.470 142.530 ;
        RECT 171.310 141.490 180.130 142.530 ;
        RECT 180.970 141.490 186.570 142.530 ;
        RECT 187.410 141.490 196.230 142.530 ;
        RECT 197.070 141.490 197.700 142.530 ;
        RECT 0.100 4.280 197.700 141.490 ;
        RECT 0.650 0.155 6.250 4.280 ;
        RECT 7.090 0.155 15.910 4.280 ;
        RECT 16.750 0.155 25.570 4.280 ;
        RECT 26.410 0.155 35.230 4.280 ;
        RECT 36.070 0.155 41.670 4.280 ;
        RECT 42.510 0.155 51.330 4.280 ;
        RECT 52.170 0.155 60.990 4.280 ;
        RECT 61.830 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 86.750 4.280 ;
        RECT 87.590 0.155 96.410 4.280 ;
        RECT 97.250 0.155 106.070 4.280 ;
        RECT 106.910 0.155 112.510 4.280 ;
        RECT 113.350 0.155 122.170 4.280 ;
        RECT 123.010 0.155 131.830 4.280 ;
        RECT 132.670 0.155 141.490 4.280 ;
        RECT 142.330 0.155 147.930 4.280 ;
        RECT 148.770 0.155 157.590 4.280 ;
        RECT 158.430 0.155 167.250 4.280 ;
        RECT 168.090 0.155 176.910 4.280 ;
        RECT 177.750 0.155 183.350 4.280 ;
        RECT 184.190 0.155 193.010 4.280 ;
        RECT 193.850 0.155 197.700 4.280 ;
      LAYER met3 ;
        RECT 4.400 139.040 197.430 139.905 ;
        RECT 4.000 130.240 197.830 139.040 ;
        RECT 4.400 128.840 197.430 130.240 ;
        RECT 4.000 123.440 197.830 128.840 ;
        RECT 4.000 122.040 197.430 123.440 ;
        RECT 4.000 120.040 197.830 122.040 ;
        RECT 4.400 118.640 197.830 120.040 ;
        RECT 4.000 113.240 197.830 118.640 ;
        RECT 4.400 111.840 197.430 113.240 ;
        RECT 4.000 103.040 197.830 111.840 ;
        RECT 4.400 101.640 197.430 103.040 ;
        RECT 4.000 92.840 197.830 101.640 ;
        RECT 4.400 91.440 197.430 92.840 ;
        RECT 4.000 86.040 197.830 91.440 ;
        RECT 4.000 84.640 197.430 86.040 ;
        RECT 4.000 82.640 197.830 84.640 ;
        RECT 4.400 81.240 197.830 82.640 ;
        RECT 4.000 75.840 197.830 81.240 ;
        RECT 4.400 74.440 197.430 75.840 ;
        RECT 4.000 65.640 197.830 74.440 ;
        RECT 4.400 64.240 197.430 65.640 ;
        RECT 4.000 55.440 197.830 64.240 ;
        RECT 4.400 54.040 197.430 55.440 ;
        RECT 4.000 48.640 197.830 54.040 ;
        RECT 4.000 47.240 197.430 48.640 ;
        RECT 4.000 45.240 197.830 47.240 ;
        RECT 4.400 43.840 197.830 45.240 ;
        RECT 4.000 38.440 197.830 43.840 ;
        RECT 4.400 37.040 197.430 38.440 ;
        RECT 4.000 28.240 197.830 37.040 ;
        RECT 4.400 26.840 197.430 28.240 ;
        RECT 4.000 18.040 197.830 26.840 ;
        RECT 4.400 16.640 197.430 18.040 ;
        RECT 4.000 11.240 197.830 16.640 ;
        RECT 4.000 9.840 197.430 11.240 ;
        RECT 4.000 7.840 197.830 9.840 ;
        RECT 4.400 6.440 197.830 7.840 ;
        RECT 4.000 1.040 197.830 6.440 ;
        RECT 4.000 0.175 197.430 1.040 ;
      LAYER met4 ;
        RECT 13.175 10.240 28.125 132.425 ;
        RECT 30.525 10.240 51.930 132.425 ;
        RECT 54.330 10.240 75.735 132.425 ;
        RECT 78.135 10.240 99.540 132.425 ;
        RECT 101.940 10.240 123.345 132.425 ;
        RECT 125.745 10.240 147.150 132.425 ;
        RECT 149.550 10.240 170.955 132.425 ;
        RECT 173.355 10.240 173.585 132.425 ;
        RECT 13.175 6.295 173.585 10.240 ;
  END
END Scalar_Register_File
END LIBRARY

