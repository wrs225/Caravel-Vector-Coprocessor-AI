magic
tech sky130A
magscale 1 2
timestamp 1692311903
<< obsli1 >>
rect 1104 2159 305532 230129
<< obsm1 >>
rect 14 892 305794 231804
<< metal2 >>
rect 18 231892 74 232692
rect 7746 231892 7802 232692
rect 16118 231892 16174 232692
rect 24490 231892 24546 232692
rect 32862 231892 32918 232692
rect 40590 231892 40646 232692
rect 48962 231892 49018 232692
rect 57334 231892 57390 232692
rect 65062 231892 65118 232692
rect 73434 231892 73490 232692
rect 81806 231892 81862 232692
rect 90178 231892 90234 232692
rect 97906 231892 97962 232692
rect 106278 231892 106334 232692
rect 114650 231892 114706 232692
rect 122378 231892 122434 232692
rect 130750 231892 130806 232692
rect 139122 231892 139178 232692
rect 147494 231892 147550 232692
rect 155222 231892 155278 232692
rect 163594 231892 163650 232692
rect 171966 231892 172022 232692
rect 179694 231892 179750 232692
rect 188066 231892 188122 232692
rect 196438 231892 196494 232692
rect 204810 231892 204866 232692
rect 212538 231892 212594 232692
rect 220910 231892 220966 232692
rect 229282 231892 229338 232692
rect 237010 231892 237066 232692
rect 245382 231892 245438 232692
rect 253754 231892 253810 232692
rect 262126 231892 262182 232692
rect 269854 231892 269910 232692
rect 278226 231892 278282 232692
rect 286598 231892 286654 232692
rect 294326 231892 294382 232692
rect 302698 231892 302754 232692
rect 18 0 74 800
rect 7746 0 7802 800
rect 16118 0 16174 800
rect 24490 0 24546 800
rect 32218 0 32274 800
rect 40590 0 40646 800
rect 48962 0 49018 800
rect 56690 0 56746 800
rect 65062 0 65118 800
rect 73434 0 73490 800
rect 81806 0 81862 800
rect 89534 0 89590 800
rect 97906 0 97962 800
rect 106278 0 106334 800
rect 114006 0 114062 800
rect 122378 0 122434 800
rect 130750 0 130806 800
rect 139122 0 139178 800
rect 146850 0 146906 800
rect 155222 0 155278 800
rect 163594 0 163650 800
rect 171322 0 171378 800
rect 179694 0 179750 800
rect 188066 0 188122 800
rect 196438 0 196494 800
rect 204166 0 204222 800
rect 212538 0 212594 800
rect 220910 0 220966 800
rect 228638 0 228694 800
rect 237010 0 237066 800
rect 245382 0 245438 800
rect 253754 0 253810 800
rect 261482 0 261538 800
rect 269854 0 269910 800
rect 278226 0 278282 800
rect 285954 0 286010 800
rect 294326 0 294382 800
rect 302698 0 302754 800
<< obsm2 >>
rect 130 231836 7690 231892
rect 7858 231836 16062 231892
rect 16230 231836 24434 231892
rect 24602 231836 32806 231892
rect 32974 231836 40534 231892
rect 40702 231836 48906 231892
rect 49074 231836 57278 231892
rect 57446 231836 65006 231892
rect 65174 231836 73378 231892
rect 73546 231836 81750 231892
rect 81918 231836 90122 231892
rect 90290 231836 97850 231892
rect 98018 231836 106222 231892
rect 106390 231836 114594 231892
rect 114762 231836 122322 231892
rect 122490 231836 130694 231892
rect 130862 231836 139066 231892
rect 139234 231836 147438 231892
rect 147606 231836 155166 231892
rect 155334 231836 163538 231892
rect 163706 231836 171910 231892
rect 172078 231836 179638 231892
rect 179806 231836 188010 231892
rect 188178 231836 196382 231892
rect 196550 231836 204754 231892
rect 204922 231836 212482 231892
rect 212650 231836 220854 231892
rect 221022 231836 229226 231892
rect 229394 231836 236954 231892
rect 237122 231836 245326 231892
rect 245494 231836 253698 231892
rect 253866 231836 262070 231892
rect 262238 231836 269798 231892
rect 269966 231836 278170 231892
rect 278338 231836 286542 231892
rect 286710 231836 294270 231892
rect 294438 231836 302642 231892
rect 302810 231836 305790 231892
rect 20 856 305790 231836
rect 130 800 7690 856
rect 7858 800 16062 856
rect 16230 800 24434 856
rect 24602 800 32162 856
rect 32330 800 40534 856
rect 40702 800 48906 856
rect 49074 800 56634 856
rect 56802 800 65006 856
rect 65174 800 73378 856
rect 73546 800 81750 856
rect 81918 800 89478 856
rect 89646 800 97850 856
rect 98018 800 106222 856
rect 106390 800 113950 856
rect 114118 800 122322 856
rect 122490 800 130694 856
rect 130862 800 139066 856
rect 139234 800 146794 856
rect 146962 800 155166 856
rect 155334 800 163538 856
rect 163706 800 171266 856
rect 171434 800 179638 856
rect 179806 800 188010 856
rect 188178 800 196382 856
rect 196550 800 204110 856
rect 204278 800 212482 856
rect 212650 800 220854 856
rect 221022 800 228582 856
rect 228750 800 236954 856
rect 237122 800 245326 856
rect 245494 800 253698 856
rect 253866 800 261426 856
rect 261594 800 269798 856
rect 269966 800 278170 856
rect 278338 800 285898 856
rect 286066 800 294270 856
rect 294438 800 302642 856
rect 302810 800 305790 856
<< metal3 >>
rect 305861 228488 306661 228608
rect 0 224408 800 224528
rect 305861 219648 306661 219768
rect 0 215568 800 215688
rect 305861 211488 306661 211608
rect 0 207408 800 207528
rect 305861 202648 306661 202768
rect 0 198568 800 198688
rect 305861 193808 306661 193928
rect 0 189728 800 189848
rect 305861 185648 306661 185768
rect 0 180888 800 181008
rect 305861 176808 306661 176928
rect 0 172728 800 172848
rect 305861 167968 306661 168088
rect 0 163888 800 164008
rect 305861 159128 306661 159248
rect 0 155048 800 155168
rect 305861 150968 306661 151088
rect 0 146888 800 147008
rect 305861 142128 306661 142248
rect 0 138048 800 138168
rect 305861 133288 306661 133408
rect 0 129208 800 129328
rect 305861 125128 306661 125248
rect 0 120368 800 120488
rect 305861 116288 306661 116408
rect 0 112208 800 112328
rect 305861 107448 306661 107568
rect 0 103368 800 103488
rect 305861 98608 306661 98728
rect 0 94528 800 94648
rect 305861 90448 306661 90568
rect 0 86368 800 86488
rect 305861 81608 306661 81728
rect 0 77528 800 77648
rect 305861 72768 306661 72888
rect 0 68688 800 68808
rect 305861 64608 306661 64728
rect 0 59848 800 59968
rect 305861 55768 306661 55888
rect 0 51688 800 51808
rect 305861 46928 306661 47048
rect 0 42848 800 42968
rect 305861 38088 306661 38208
rect 0 34008 800 34128
rect 305861 29928 306661 30048
rect 0 25848 800 25968
rect 305861 21088 306661 21208
rect 0 17008 800 17128
rect 305861 12248 306661 12368
rect 0 8168 800 8288
rect 305861 4088 306661 4208
<< obsm3 >>
rect 800 228688 305861 230349
rect 800 228408 305781 228688
rect 800 224608 305861 228408
rect 880 224328 305861 224608
rect 800 219848 305861 224328
rect 800 219568 305781 219848
rect 800 215768 305861 219568
rect 880 215488 305861 215768
rect 800 211688 305861 215488
rect 800 211408 305781 211688
rect 800 207608 305861 211408
rect 880 207328 305861 207608
rect 800 202848 305861 207328
rect 800 202568 305781 202848
rect 800 198768 305861 202568
rect 880 198488 305861 198768
rect 800 194008 305861 198488
rect 800 193728 305781 194008
rect 800 189928 305861 193728
rect 880 189648 305861 189928
rect 800 185848 305861 189648
rect 800 185568 305781 185848
rect 800 181088 305861 185568
rect 880 180808 305861 181088
rect 800 177008 305861 180808
rect 800 176728 305781 177008
rect 800 172928 305861 176728
rect 880 172648 305861 172928
rect 800 168168 305861 172648
rect 800 167888 305781 168168
rect 800 164088 305861 167888
rect 880 163808 305861 164088
rect 800 159328 305861 163808
rect 800 159048 305781 159328
rect 800 155248 305861 159048
rect 880 154968 305861 155248
rect 800 151168 305861 154968
rect 800 150888 305781 151168
rect 800 147088 305861 150888
rect 880 146808 305861 147088
rect 800 142328 305861 146808
rect 800 142048 305781 142328
rect 800 138248 305861 142048
rect 880 137968 305861 138248
rect 800 133488 305861 137968
rect 800 133208 305781 133488
rect 800 129408 305861 133208
rect 880 129128 305861 129408
rect 800 125328 305861 129128
rect 800 125048 305781 125328
rect 800 120568 305861 125048
rect 880 120288 305861 120568
rect 800 116488 305861 120288
rect 800 116208 305781 116488
rect 800 112408 305861 116208
rect 880 112128 305861 112408
rect 800 107648 305861 112128
rect 800 107368 305781 107648
rect 800 103568 305861 107368
rect 880 103288 305861 103568
rect 800 98808 305861 103288
rect 800 98528 305781 98808
rect 800 94728 305861 98528
rect 880 94448 305861 94728
rect 800 90648 305861 94448
rect 800 90368 305781 90648
rect 800 86568 305861 90368
rect 880 86288 305861 86568
rect 800 81808 305861 86288
rect 800 81528 305781 81808
rect 800 77728 305861 81528
rect 880 77448 305861 77728
rect 800 72968 305861 77448
rect 800 72688 305781 72968
rect 800 68888 305861 72688
rect 880 68608 305861 68888
rect 800 64808 305861 68608
rect 800 64528 305781 64808
rect 800 60048 305861 64528
rect 880 59768 305861 60048
rect 800 55968 305861 59768
rect 800 55688 305781 55968
rect 800 51888 305861 55688
rect 880 51608 305861 51888
rect 800 47128 305861 51608
rect 800 46848 305781 47128
rect 800 43048 305861 46848
rect 880 42768 305861 43048
rect 800 38288 305861 42768
rect 800 38008 305781 38288
rect 800 34208 305861 38008
rect 880 33928 305861 34208
rect 800 30128 305861 33928
rect 800 29848 305781 30128
rect 800 26048 305861 29848
rect 880 25768 305861 26048
rect 800 21288 305861 25768
rect 800 21008 305781 21288
rect 800 17208 305861 21008
rect 880 16928 305861 17208
rect 800 12448 305861 16928
rect 800 12168 305781 12448
rect 800 8368 305861 12168
rect 880 8088 305861 8368
rect 800 4288 305861 8088
rect 800 4008 305781 4288
rect 800 1803 305861 4008
<< metal4 >>
rect 4208 2128 4528 230160
rect 19568 2128 19888 230160
rect 34928 2128 35248 230160
rect 50288 2128 50608 230160
rect 65648 2128 65968 230160
rect 81008 2128 81328 230160
rect 96368 2128 96688 230160
rect 111728 2128 112048 230160
rect 127088 2128 127408 230160
rect 142448 2128 142768 230160
rect 157808 2128 158128 230160
rect 173168 2128 173488 230160
rect 188528 2128 188848 230160
rect 203888 2128 204208 230160
rect 219248 2128 219568 230160
rect 234608 2128 234928 230160
rect 249968 2128 250288 230160
rect 265328 2128 265648 230160
rect 280688 2128 281008 230160
rect 296048 2128 296368 230160
<< obsm4 >>
rect 7235 230240 289189 230349
rect 7235 2048 19488 230240
rect 19968 2048 34848 230240
rect 35328 2048 50208 230240
rect 50688 2048 65568 230240
rect 66048 2048 80928 230240
rect 81408 2048 96288 230240
rect 96768 2048 111648 230240
rect 112128 2048 127008 230240
rect 127488 2048 142368 230240
rect 142848 2048 157728 230240
rect 158208 2048 173088 230240
rect 173568 2048 188448 230240
rect 188928 2048 203808 230240
rect 204288 2048 219168 230240
rect 219648 2048 234528 230240
rect 235008 2048 249888 230240
rect 250368 2048 265248 230240
rect 265728 2048 280608 230240
rect 281088 2048 289189 230240
rect 7235 1803 289189 2048
<< labels >>
rlabel metal2 s 18 231892 74 232692 6 clk
port 1 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 rAddr1_1[0]
port 2 nsew signal input
rlabel metal3 s 0 189728 800 189848 6 rAddr1_1[1]
port 3 nsew signal input
rlabel metal2 s 155222 231892 155278 232692 6 rAddr1_1[2]
port 4 nsew signal input
rlabel metal3 s 305861 228488 306661 228608 6 rAddr1_1[3]
port 5 nsew signal input
rlabel metal3 s 0 215568 800 215688 6 rAddr1_1[4]
port 6 nsew signal input
rlabel metal2 s 278226 231892 278282 232692 6 rAddr1_2[0]
port 7 nsew signal input
rlabel metal2 s 253754 0 253810 800 6 rAddr1_2[1]
port 8 nsew signal input
rlabel metal2 s 81806 231892 81862 232692 6 rAddr1_2[2]
port 9 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 rAddr1_2[3]
port 10 nsew signal input
rlabel metal2 s 262126 231892 262182 232692 6 rAddr1_2[4]
port 11 nsew signal input
rlabel metal3 s 305861 64608 306661 64728 6 rAddr2_1[0]
port 12 nsew signal input
rlabel metal2 s 269854 231892 269910 232692 6 rAddr2_1[1]
port 13 nsew signal input
rlabel metal3 s 0 163888 800 164008 6 rAddr2_1[2]
port 14 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 rAddr2_1[3]
port 15 nsew signal input
rlabel metal2 s 147494 231892 147550 232692 6 rAddr2_1[4]
port 16 nsew signal input
rlabel metal3 s 305861 55768 306661 55888 6 rAddr2_2[0]
port 17 nsew signal input
rlabel metal2 s 163594 231892 163650 232692 6 rAddr2_2[1]
port 18 nsew signal input
rlabel metal3 s 305861 159128 306661 159248 6 rAddr2_2[2]
port 19 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 rAddr2_2[3]
port 20 nsew signal input
rlabel metal3 s 305861 116288 306661 116408 6 rAddr2_2[4]
port 21 nsew signal input
rlabel metal3 s 305861 107448 306661 107568 6 rData1[0]
port 22 nsew signal output
rlabel metal2 s 97906 231892 97962 232692 6 rData1[10]
port 23 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 rData1[11]
port 24 nsew signal output
rlabel metal2 s 220910 0 220966 800 6 rData1[12]
port 25 nsew signal output
rlabel metal3 s 305861 125128 306661 125248 6 rData1[13]
port 26 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 rData1[14]
port 27 nsew signal output
rlabel metal3 s 0 146888 800 147008 6 rData1[15]
port 28 nsew signal output
rlabel metal2 s 302698 0 302754 800 6 rData1[16]
port 29 nsew signal output
rlabel metal3 s 305861 150968 306661 151088 6 rData1[17]
port 30 nsew signal output
rlabel metal2 s 204810 231892 204866 232692 6 rData1[18]
port 31 nsew signal output
rlabel metal2 s 261482 0 261538 800 6 rData1[19]
port 32 nsew signal output
rlabel metal2 s 65062 231892 65118 232692 6 rData1[1]
port 33 nsew signal output
rlabel metal3 s 305861 38088 306661 38208 6 rData1[20]
port 34 nsew signal output
rlabel metal2 s 32862 231892 32918 232692 6 rData1[21]
port 35 nsew signal output
rlabel metal3 s 0 207408 800 207528 6 rData1[22]
port 36 nsew signal output
rlabel metal2 s 294326 231892 294382 232692 6 rData1[23]
port 37 nsew signal output
rlabel metal2 s 228638 0 228694 800 6 rData1[24]
port 38 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 rData1[25]
port 39 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 rData1[26]
port 40 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 rData1[27]
port 41 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 rData1[28]
port 42 nsew signal output
rlabel metal3 s 305861 12248 306661 12368 6 rData1[29]
port 43 nsew signal output
rlabel metal2 s 188066 231892 188122 232692 6 rData1[2]
port 44 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 rData1[30]
port 45 nsew signal output
rlabel metal2 s 229282 231892 229338 232692 6 rData1[31]
port 46 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 rData1[3]
port 47 nsew signal output
rlabel metal2 s 302698 231892 302754 232692 6 rData1[4]
port 48 nsew signal output
rlabel metal2 s 114650 231892 114706 232692 6 rData1[5]
port 49 nsew signal output
rlabel metal2 s 278226 0 278282 800 6 rData1[6]
port 50 nsew signal output
rlabel metal3 s 305861 167968 306661 168088 6 rData1[7]
port 51 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 rData1[8]
port 52 nsew signal output
rlabel metal2 s 179694 231892 179750 232692 6 rData1[9]
port 53 nsew signal output
rlabel metal2 s 130750 231892 130806 232692 6 rData2[0]
port 54 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 rData2[10]
port 55 nsew signal output
rlabel metal3 s 305861 219648 306661 219768 6 rData2[11]
port 56 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 rData2[12]
port 57 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 rData2[13]
port 58 nsew signal output
rlabel metal2 s 106278 231892 106334 232692 6 rData2[14]
port 59 nsew signal output
rlabel metal3 s 0 172728 800 172848 6 rData2[15]
port 60 nsew signal output
rlabel metal3 s 305861 202648 306661 202768 6 rData2[16]
port 61 nsew signal output
rlabel metal2 s 57334 231892 57390 232692 6 rData2[17]
port 62 nsew signal output
rlabel metal3 s 305861 185648 306661 185768 6 rData2[18]
port 63 nsew signal output
rlabel metal2 s 73434 231892 73490 232692 6 rData2[19]
port 64 nsew signal output
rlabel metal2 s 139122 231892 139178 232692 6 rData2[1]
port 65 nsew signal output
rlabel metal2 s 220910 231892 220966 232692 6 rData2[20]
port 66 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 rData2[21]
port 67 nsew signal output
rlabel metal3 s 305861 72768 306661 72888 6 rData2[22]
port 68 nsew signal output
rlabel metal3 s 305861 29928 306661 30048 6 rData2[23]
port 69 nsew signal output
rlabel metal3 s 0 198568 800 198688 6 rData2[24]
port 70 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 rData2[25]
port 71 nsew signal output
rlabel metal2 s 269854 0 269910 800 6 rData2[26]
port 72 nsew signal output
rlabel metal3 s 305861 46928 306661 47048 6 rData2[27]
port 73 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 rData2[28]
port 74 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 rData2[29]
port 75 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 rData2[2]
port 76 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 rData2[30]
port 77 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 rData2[31]
port 78 nsew signal output
rlabel metal3 s 305861 211488 306661 211608 6 rData2[3]
port 79 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 rData2[4]
port 80 nsew signal output
rlabel metal2 s 294326 0 294382 800 6 rData2[5]
port 81 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 rData2[6]
port 82 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 rData2[7]
port 83 nsew signal output
rlabel metal2 s 171966 231892 172022 232692 6 rData2[8]
port 84 nsew signal output
rlabel metal2 s 196438 0 196494 800 6 rData2[9]
port 85 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 reset
port 86 nsew signal input
rlabel metal4 s 4208 2128 4528 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 230160 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 230160 6 vssd1
port 88 nsew ground bidirectional
rlabel metal2 s 97906 0 97962 800 6 wAddr1[0]
port 89 nsew signal input
rlabel metal2 s 285954 0 286010 800 6 wAddr1[1]
port 90 nsew signal input
rlabel metal3 s 305861 142128 306661 142248 6 wAddr1[2]
port 91 nsew signal input
rlabel metal3 s 305861 81608 306661 81728 6 wAddr1[3]
port 92 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 wAddr1[4]
port 93 nsew signal input
rlabel metal3 s 0 180888 800 181008 6 wAddr2[0]
port 94 nsew signal input
rlabel metal3 s 305861 21088 306661 21208 6 wAddr2[1]
port 95 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wAddr2[2]
port 96 nsew signal input
rlabel metal3 s 305861 98608 306661 98728 6 wAddr2[3]
port 97 nsew signal input
rlabel metal3 s 305861 176808 306661 176928 6 wAddr2[4]
port 98 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 wData[0]
port 99 nsew signal input
rlabel metal3 s 305861 193808 306661 193928 6 wData[10]
port 100 nsew signal input
rlabel metal2 s 16118 231892 16174 232692 6 wData[11]
port 101 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 wData[12]
port 102 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 wData[13]
port 103 nsew signal input
rlabel metal2 s 18 0 74 800 6 wData[14]
port 104 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 wData[15]
port 105 nsew signal input
rlabel metal2 s 40590 231892 40646 232692 6 wData[16]
port 106 nsew signal input
rlabel metal2 s 122378 231892 122434 232692 6 wData[17]
port 107 nsew signal input
rlabel metal2 s 212538 231892 212594 232692 6 wData[18]
port 108 nsew signal input
rlabel metal3 s 0 224408 800 224528 6 wData[19]
port 109 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 wData[1]
port 110 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wData[20]
port 111 nsew signal input
rlabel metal2 s 253754 231892 253810 232692 6 wData[21]
port 112 nsew signal input
rlabel metal2 s 196438 231892 196494 232692 6 wData[22]
port 113 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 wData[23]
port 114 nsew signal input
rlabel metal2 s 286598 231892 286654 232692 6 wData[24]
port 115 nsew signal input
rlabel metal3 s 305861 4088 306661 4208 6 wData[25]
port 116 nsew signal input
rlabel metal2 s 24490 231892 24546 232692 6 wData[26]
port 117 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 wData[27]
port 118 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wData[28]
port 119 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 wData[29]
port 120 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wData[2]
port 121 nsew signal input
rlabel metal3 s 305861 133288 306661 133408 6 wData[30]
port 122 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 wData[31]
port 123 nsew signal input
rlabel metal2 s 245382 231892 245438 232692 6 wData[3]
port 124 nsew signal input
rlabel metal2 s 237010 231892 237066 232692 6 wData[4]
port 125 nsew signal input
rlabel metal2 s 48962 231892 49018 232692 6 wData[5]
port 126 nsew signal input
rlabel metal2 s 90178 231892 90234 232692 6 wData[6]
port 127 nsew signal input
rlabel metal2 s 188066 0 188122 800 6 wData[7]
port 128 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wData[8]
port 129 nsew signal input
rlabel metal2 s 7746 231892 7802 232692 6 wData[9]
port 130 nsew signal input
rlabel metal3 s 305861 90448 306661 90568 6 wEnable
port 131 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 306661 232692
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 123636628
string GDS_FILE /home/courtney/Desktop/Caravel-Vector-Coprocessor-AI/openlane/VectorRegFile/runs/23_08_17_17_16/results/signoff/VectorRegFile.magic.gds
string GDS_START 657464
<< end >>

