VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO VectorRegFile
  CLASS BLOCK ;
  FOREIGN VectorRegFile ;
  ORIGIN 0.000 0.000 ;
  SIZE 1533.305 BY 1163.460 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1159.460 0.370 1163.460 ;
    END
  END clk
  PIN rAddr1_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END rAddr1_1[0]
  PIN rAddr1_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END rAddr1_1[1]
  PIN rAddr1_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 1159.460 776.390 1163.460 ;
    END
  END rAddr1_1[2]
  PIN rAddr1_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 1142.440 1533.305 1143.040 ;
    END
  END rAddr1_1[3]
  PIN rAddr1_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END rAddr1_1[4]
  PIN rAddr1_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 1159.460 1391.410 1163.460 ;
    END
  END rAddr1_2[0]
  PIN rAddr1_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 4.000 ;
    END
  END rAddr1_2[1]
  PIN rAddr1_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 1159.460 409.310 1163.460 ;
    END
  END rAddr1_2[2]
  PIN rAddr1_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END rAddr1_2[3]
  PIN rAddr1_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 1159.460 1310.910 1163.460 ;
    END
  END rAddr1_2[4]
  PIN rAddr2_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 323.040 1533.305 323.640 ;
    END
  END rAddr2_1[0]
  PIN rAddr2_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 1159.460 1349.550 1163.460 ;
    END
  END rAddr2_1[1]
  PIN rAddr2_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END rAddr2_1[2]
  PIN rAddr2_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END rAddr2_1[3]
  PIN rAddr2_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 1159.460 737.750 1163.460 ;
    END
  END rAddr2_1[4]
  PIN rAddr2_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 278.840 1533.305 279.440 ;
    END
  END rAddr2_2[0]
  PIN rAddr2_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 1159.460 818.250 1163.460 ;
    END
  END rAddr2_2[1]
  PIN rAddr2_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 795.640 1533.305 796.240 ;
    END
  END rAddr2_2[2]
  PIN rAddr2_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END rAddr2_2[3]
  PIN rAddr2_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 581.440 1533.305 582.040 ;
    END
  END rAddr2_2[4]
  PIN rData1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 537.240 1533.305 537.840 ;
    END
  END rData1[0]
  PIN rData1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 1159.460 489.810 1163.460 ;
    END
  END rData1[10]
  PIN rData1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END rData1[11]
  PIN rData1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END rData1[12]
  PIN rData1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 625.640 1533.305 626.240 ;
    END
  END rData1[13]
  PIN rData1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END rData1[14]
  PIN rData1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END rData1[15]
  PIN rData1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 0.000 1513.770 4.000 ;
    END
  END rData1[16]
  PIN rData1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 754.840 1533.305 755.440 ;
    END
  END rData1[17]
  PIN rData1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 1159.460 1024.330 1163.460 ;
    END
  END rData1[18]
  PIN rData1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END rData1[19]
  PIN rData1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 1159.460 325.590 1163.460 ;
    END
  END rData1[1]
  PIN rData1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 190.440 1533.305 191.040 ;
    END
  END rData1[20]
  PIN rData1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 1159.460 164.590 1163.460 ;
    END
  END rData1[21]
  PIN rData1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END rData1[22]
  PIN rData1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 1159.460 1471.910 1163.460 ;
    END
  END rData1[23]
  PIN rData1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END rData1[24]
  PIN rData1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END rData1[25]
  PIN rData1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END rData1[26]
  PIN rData1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END rData1[27]
  PIN rData1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END rData1[28]
  PIN rData1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 61.240 1533.305 61.840 ;
    END
  END rData1[29]
  PIN rData1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 1159.460 940.610 1163.460 ;
    END
  END rData1[2]
  PIN rData1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END rData1[30]
  PIN rData1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 1159.460 1146.690 1163.460 ;
    END
  END rData1[31]
  PIN rData1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END rData1[3]
  PIN rData1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 1159.460 1513.770 1163.460 ;
    END
  END rData1[4]
  PIN rData1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 1159.460 573.530 1163.460 ;
    END
  END rData1[5]
  PIN rData1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END rData1[6]
  PIN rData1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 839.840 1533.305 840.440 ;
    END
  END rData1[7]
  PIN rData1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END rData1[8]
  PIN rData1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 1159.460 898.750 1163.460 ;
    END
  END rData1[9]
  PIN rData2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1159.460 654.030 1163.460 ;
    END
  END rData2[0]
  PIN rData2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END rData2[10]
  PIN rData2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 1098.240 1533.305 1098.840 ;
    END
  END rData2[11]
  PIN rData2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END rData2[12]
  PIN rData2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END rData2[13]
  PIN rData2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 1159.460 531.670 1163.460 ;
    END
  END rData2[14]
  PIN rData2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END rData2[15]
  PIN rData2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 1013.240 1533.305 1013.840 ;
    END
  END rData2[16]
  PIN rData2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 1159.460 286.950 1163.460 ;
    END
  END rData2[17]
  PIN rData2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 928.240 1533.305 928.840 ;
    END
  END rData2[18]
  PIN rData2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 1159.460 367.450 1163.460 ;
    END
  END rData2[19]
  PIN rData2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 1159.460 695.890 1163.460 ;
    END
  END rData2[1]
  PIN rData2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 1159.460 1104.830 1163.460 ;
    END
  END rData2[20]
  PIN rData2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END rData2[21]
  PIN rData2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 363.840 1533.305 364.440 ;
    END
  END rData2[22]
  PIN rData2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 149.640 1533.305 150.240 ;
    END
  END rData2[23]
  PIN rData2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END rData2[24]
  PIN rData2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END rData2[25]
  PIN rData2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END rData2[26]
  PIN rData2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 234.640 1533.305 235.240 ;
    END
  END rData2[27]
  PIN rData2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END rData2[28]
  PIN rData2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END rData2[29]
  PIN rData2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END rData2[2]
  PIN rData2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END rData2[30]
  PIN rData2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END rData2[31]
  PIN rData2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 1057.440 1533.305 1058.040 ;
    END
  END rData2[3]
  PIN rData2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END rData2[4]
  PIN rData2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 4.000 ;
    END
  END rData2[5]
  PIN rData2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END rData2[6]
  PIN rData2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END rData2[7]
  PIN rData2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 1159.460 860.110 1163.460 ;
    END
  END rData2[8]
  PIN rData2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END rData2[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1150.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1150.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1150.800 ;
    END
  END vssd1
  PIN wAddr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END wAddr1[0]
  PIN wAddr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END wAddr1[1]
  PIN wAddr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 710.640 1533.305 711.240 ;
    END
  END wAddr1[2]
  PIN wAddr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 408.040 1533.305 408.640 ;
    END
  END wAddr1[3]
  PIN wAddr1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END wAddr1[4]
  PIN wAddr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END wAddr2[0]
  PIN wAddr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 105.440 1533.305 106.040 ;
    END
  END wAddr2[1]
  PIN wAddr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END wAddr2[2]
  PIN wAddr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 493.040 1533.305 493.640 ;
    END
  END wAddr2[3]
  PIN wAddr2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 884.040 1533.305 884.640 ;
    END
  END wAddr2[4]
  PIN wData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 0.000 1185.330 4.000 ;
    END
  END wData[0]
  PIN wData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 969.040 1533.305 969.640 ;
    END
  END wData[10]
  PIN wData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1159.460 80.870 1163.460 ;
    END
  END wData[11]
  PIN wData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END wData[12]
  PIN wData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END wData[13]
  PIN wData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wData[14]
  PIN wData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END wData[15]
  PIN wData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 1159.460 203.230 1163.460 ;
    END
  END wData[16]
  PIN wData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1159.460 612.170 1163.460 ;
    END
  END wData[17]
  PIN wData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 1159.460 1062.970 1163.460 ;
    END
  END wData[18]
  PIN wData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END wData[19]
  PIN wData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END wData[1]
  PIN wData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wData[20]
  PIN wData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 1159.460 1269.050 1163.460 ;
    END
  END wData[21]
  PIN wData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 1159.460 982.470 1163.460 ;
    END
  END wData[22]
  PIN wData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END wData[23]
  PIN wData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 1159.460 1433.270 1163.460 ;
    END
  END wData[24]
  PIN wData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 20.440 1533.305 21.040 ;
    END
  END wData[25]
  PIN wData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1159.460 122.730 1163.460 ;
    END
  END wData[26]
  PIN wData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END wData[27]
  PIN wData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wData[28]
  PIN wData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END wData[29]
  PIN wData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wData[2]
  PIN wData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 666.440 1533.305 667.040 ;
    END
  END wData[30]
  PIN wData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END wData[31]
  PIN wData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 1159.460 1227.190 1163.460 ;
    END
  END wData[3]
  PIN wData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 1159.460 1185.330 1163.460 ;
    END
  END wData[4]
  PIN wData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 1159.460 245.090 1163.460 ;
    END
  END wData[5]
  PIN wData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 1159.460 451.170 1163.460 ;
    END
  END wData[6]
  PIN wData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END wData[7]
  PIN wData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END wData[8]
  PIN wData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1159.460 39.010 1163.460 ;
    END
  END wData[9]
  PIN wEnable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.305 452.240 1533.305 452.840 ;
    END
  END wEnable
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1527.660 1150.645 ;
      LAYER met1 ;
        RECT 0.070 4.460 1528.970 1159.020 ;
      LAYER met2 ;
        RECT 0.650 1159.180 38.450 1159.460 ;
        RECT 39.290 1159.180 80.310 1159.460 ;
        RECT 81.150 1159.180 122.170 1159.460 ;
        RECT 123.010 1159.180 164.030 1159.460 ;
        RECT 164.870 1159.180 202.670 1159.460 ;
        RECT 203.510 1159.180 244.530 1159.460 ;
        RECT 245.370 1159.180 286.390 1159.460 ;
        RECT 287.230 1159.180 325.030 1159.460 ;
        RECT 325.870 1159.180 366.890 1159.460 ;
        RECT 367.730 1159.180 408.750 1159.460 ;
        RECT 409.590 1159.180 450.610 1159.460 ;
        RECT 451.450 1159.180 489.250 1159.460 ;
        RECT 490.090 1159.180 531.110 1159.460 ;
        RECT 531.950 1159.180 572.970 1159.460 ;
        RECT 573.810 1159.180 611.610 1159.460 ;
        RECT 612.450 1159.180 653.470 1159.460 ;
        RECT 654.310 1159.180 695.330 1159.460 ;
        RECT 696.170 1159.180 737.190 1159.460 ;
        RECT 738.030 1159.180 775.830 1159.460 ;
        RECT 776.670 1159.180 817.690 1159.460 ;
        RECT 818.530 1159.180 859.550 1159.460 ;
        RECT 860.390 1159.180 898.190 1159.460 ;
        RECT 899.030 1159.180 940.050 1159.460 ;
        RECT 940.890 1159.180 981.910 1159.460 ;
        RECT 982.750 1159.180 1023.770 1159.460 ;
        RECT 1024.610 1159.180 1062.410 1159.460 ;
        RECT 1063.250 1159.180 1104.270 1159.460 ;
        RECT 1105.110 1159.180 1146.130 1159.460 ;
        RECT 1146.970 1159.180 1184.770 1159.460 ;
        RECT 1185.610 1159.180 1226.630 1159.460 ;
        RECT 1227.470 1159.180 1268.490 1159.460 ;
        RECT 1269.330 1159.180 1310.350 1159.460 ;
        RECT 1311.190 1159.180 1348.990 1159.460 ;
        RECT 1349.830 1159.180 1390.850 1159.460 ;
        RECT 1391.690 1159.180 1432.710 1159.460 ;
        RECT 1433.550 1159.180 1471.350 1159.460 ;
        RECT 1472.190 1159.180 1513.210 1159.460 ;
        RECT 1514.050 1159.180 1528.950 1159.460 ;
        RECT 0.100 4.280 1528.950 1159.180 ;
        RECT 0.650 4.000 38.450 4.280 ;
        RECT 39.290 4.000 80.310 4.280 ;
        RECT 81.150 4.000 122.170 4.280 ;
        RECT 123.010 4.000 160.810 4.280 ;
        RECT 161.650 4.000 202.670 4.280 ;
        RECT 203.510 4.000 244.530 4.280 ;
        RECT 245.370 4.000 283.170 4.280 ;
        RECT 284.010 4.000 325.030 4.280 ;
        RECT 325.870 4.000 366.890 4.280 ;
        RECT 367.730 4.000 408.750 4.280 ;
        RECT 409.590 4.000 447.390 4.280 ;
        RECT 448.230 4.000 489.250 4.280 ;
        RECT 490.090 4.000 531.110 4.280 ;
        RECT 531.950 4.000 569.750 4.280 ;
        RECT 570.590 4.000 611.610 4.280 ;
        RECT 612.450 4.000 653.470 4.280 ;
        RECT 654.310 4.000 695.330 4.280 ;
        RECT 696.170 4.000 733.970 4.280 ;
        RECT 734.810 4.000 775.830 4.280 ;
        RECT 776.670 4.000 817.690 4.280 ;
        RECT 818.530 4.000 856.330 4.280 ;
        RECT 857.170 4.000 898.190 4.280 ;
        RECT 899.030 4.000 940.050 4.280 ;
        RECT 940.890 4.000 981.910 4.280 ;
        RECT 982.750 4.000 1020.550 4.280 ;
        RECT 1021.390 4.000 1062.410 4.280 ;
        RECT 1063.250 4.000 1104.270 4.280 ;
        RECT 1105.110 4.000 1142.910 4.280 ;
        RECT 1143.750 4.000 1184.770 4.280 ;
        RECT 1185.610 4.000 1226.630 4.280 ;
        RECT 1227.470 4.000 1268.490 4.280 ;
        RECT 1269.330 4.000 1307.130 4.280 ;
        RECT 1307.970 4.000 1348.990 4.280 ;
        RECT 1349.830 4.000 1390.850 4.280 ;
        RECT 1391.690 4.000 1429.490 4.280 ;
        RECT 1430.330 4.000 1471.350 4.280 ;
        RECT 1472.190 4.000 1513.210 4.280 ;
        RECT 1514.050 4.000 1528.950 4.280 ;
      LAYER met3 ;
        RECT 4.000 1143.440 1529.305 1151.745 ;
        RECT 4.000 1142.040 1528.905 1143.440 ;
        RECT 4.000 1123.040 1529.305 1142.040 ;
        RECT 4.400 1121.640 1529.305 1123.040 ;
        RECT 4.000 1099.240 1529.305 1121.640 ;
        RECT 4.000 1097.840 1528.905 1099.240 ;
        RECT 4.000 1078.840 1529.305 1097.840 ;
        RECT 4.400 1077.440 1529.305 1078.840 ;
        RECT 4.000 1058.440 1529.305 1077.440 ;
        RECT 4.000 1057.040 1528.905 1058.440 ;
        RECT 4.000 1038.040 1529.305 1057.040 ;
        RECT 4.400 1036.640 1529.305 1038.040 ;
        RECT 4.000 1014.240 1529.305 1036.640 ;
        RECT 4.000 1012.840 1528.905 1014.240 ;
        RECT 4.000 993.840 1529.305 1012.840 ;
        RECT 4.400 992.440 1529.305 993.840 ;
        RECT 4.000 970.040 1529.305 992.440 ;
        RECT 4.000 968.640 1528.905 970.040 ;
        RECT 4.000 949.640 1529.305 968.640 ;
        RECT 4.400 948.240 1529.305 949.640 ;
        RECT 4.000 929.240 1529.305 948.240 ;
        RECT 4.000 927.840 1528.905 929.240 ;
        RECT 4.000 905.440 1529.305 927.840 ;
        RECT 4.400 904.040 1529.305 905.440 ;
        RECT 4.000 885.040 1529.305 904.040 ;
        RECT 4.000 883.640 1528.905 885.040 ;
        RECT 4.000 864.640 1529.305 883.640 ;
        RECT 4.400 863.240 1529.305 864.640 ;
        RECT 4.000 840.840 1529.305 863.240 ;
        RECT 4.000 839.440 1528.905 840.840 ;
        RECT 4.000 820.440 1529.305 839.440 ;
        RECT 4.400 819.040 1529.305 820.440 ;
        RECT 4.000 796.640 1529.305 819.040 ;
        RECT 4.000 795.240 1528.905 796.640 ;
        RECT 4.000 776.240 1529.305 795.240 ;
        RECT 4.400 774.840 1529.305 776.240 ;
        RECT 4.000 755.840 1529.305 774.840 ;
        RECT 4.000 754.440 1528.905 755.840 ;
        RECT 4.000 735.440 1529.305 754.440 ;
        RECT 4.400 734.040 1529.305 735.440 ;
        RECT 4.000 711.640 1529.305 734.040 ;
        RECT 4.000 710.240 1528.905 711.640 ;
        RECT 4.000 691.240 1529.305 710.240 ;
        RECT 4.400 689.840 1529.305 691.240 ;
        RECT 4.000 667.440 1529.305 689.840 ;
        RECT 4.000 666.040 1528.905 667.440 ;
        RECT 4.000 647.040 1529.305 666.040 ;
        RECT 4.400 645.640 1529.305 647.040 ;
        RECT 4.000 626.640 1529.305 645.640 ;
        RECT 4.000 625.240 1528.905 626.640 ;
        RECT 4.000 602.840 1529.305 625.240 ;
        RECT 4.400 601.440 1529.305 602.840 ;
        RECT 4.000 582.440 1529.305 601.440 ;
        RECT 4.000 581.040 1528.905 582.440 ;
        RECT 4.000 562.040 1529.305 581.040 ;
        RECT 4.400 560.640 1529.305 562.040 ;
        RECT 4.000 538.240 1529.305 560.640 ;
        RECT 4.000 536.840 1528.905 538.240 ;
        RECT 4.000 517.840 1529.305 536.840 ;
        RECT 4.400 516.440 1529.305 517.840 ;
        RECT 4.000 494.040 1529.305 516.440 ;
        RECT 4.000 492.640 1528.905 494.040 ;
        RECT 4.000 473.640 1529.305 492.640 ;
        RECT 4.400 472.240 1529.305 473.640 ;
        RECT 4.000 453.240 1529.305 472.240 ;
        RECT 4.000 451.840 1528.905 453.240 ;
        RECT 4.000 432.840 1529.305 451.840 ;
        RECT 4.400 431.440 1529.305 432.840 ;
        RECT 4.000 409.040 1529.305 431.440 ;
        RECT 4.000 407.640 1528.905 409.040 ;
        RECT 4.000 388.640 1529.305 407.640 ;
        RECT 4.400 387.240 1529.305 388.640 ;
        RECT 4.000 364.840 1529.305 387.240 ;
        RECT 4.000 363.440 1528.905 364.840 ;
        RECT 4.000 344.440 1529.305 363.440 ;
        RECT 4.400 343.040 1529.305 344.440 ;
        RECT 4.000 324.040 1529.305 343.040 ;
        RECT 4.000 322.640 1528.905 324.040 ;
        RECT 4.000 300.240 1529.305 322.640 ;
        RECT 4.400 298.840 1529.305 300.240 ;
        RECT 4.000 279.840 1529.305 298.840 ;
        RECT 4.000 278.440 1528.905 279.840 ;
        RECT 4.000 259.440 1529.305 278.440 ;
        RECT 4.400 258.040 1529.305 259.440 ;
        RECT 4.000 235.640 1529.305 258.040 ;
        RECT 4.000 234.240 1528.905 235.640 ;
        RECT 4.000 215.240 1529.305 234.240 ;
        RECT 4.400 213.840 1529.305 215.240 ;
        RECT 4.000 191.440 1529.305 213.840 ;
        RECT 4.000 190.040 1528.905 191.440 ;
        RECT 4.000 171.040 1529.305 190.040 ;
        RECT 4.400 169.640 1529.305 171.040 ;
        RECT 4.000 150.640 1529.305 169.640 ;
        RECT 4.000 149.240 1528.905 150.640 ;
        RECT 4.000 130.240 1529.305 149.240 ;
        RECT 4.400 128.840 1529.305 130.240 ;
        RECT 4.000 106.440 1529.305 128.840 ;
        RECT 4.000 105.040 1528.905 106.440 ;
        RECT 4.000 86.040 1529.305 105.040 ;
        RECT 4.400 84.640 1529.305 86.040 ;
        RECT 4.000 62.240 1529.305 84.640 ;
        RECT 4.000 60.840 1528.905 62.240 ;
        RECT 4.000 41.840 1529.305 60.840 ;
        RECT 4.400 40.440 1529.305 41.840 ;
        RECT 4.000 21.440 1529.305 40.440 ;
        RECT 4.000 20.040 1528.905 21.440 ;
        RECT 4.000 9.015 1529.305 20.040 ;
      LAYER met4 ;
        RECT 36.175 1151.200 1445.945 1151.745 ;
        RECT 36.175 10.240 97.440 1151.200 ;
        RECT 99.840 10.240 174.240 1151.200 ;
        RECT 176.640 10.240 251.040 1151.200 ;
        RECT 253.440 10.240 327.840 1151.200 ;
        RECT 330.240 10.240 404.640 1151.200 ;
        RECT 407.040 10.240 481.440 1151.200 ;
        RECT 483.840 10.240 558.240 1151.200 ;
        RECT 560.640 10.240 635.040 1151.200 ;
        RECT 637.440 10.240 711.840 1151.200 ;
        RECT 714.240 10.240 788.640 1151.200 ;
        RECT 791.040 10.240 865.440 1151.200 ;
        RECT 867.840 10.240 942.240 1151.200 ;
        RECT 944.640 10.240 1019.040 1151.200 ;
        RECT 1021.440 10.240 1095.840 1151.200 ;
        RECT 1098.240 10.240 1172.640 1151.200 ;
        RECT 1175.040 10.240 1249.440 1151.200 ;
        RECT 1251.840 10.240 1326.240 1151.200 ;
        RECT 1328.640 10.240 1403.040 1151.200 ;
        RECT 1405.440 10.240 1445.945 1151.200 ;
        RECT 36.175 9.015 1445.945 10.240 ;
  END
END VectorRegFile
END LIBRARY

